      if(sum_current[i] == sum_value && co_current[i] == co_value) begin
        fitness[i] = fitness[i] + 1;
      end
