input logic clk
input logic rst
input logic i
output logic out
