`timescale 1ps/1ps
// Include all individivuals
`include "tmp/individual_0.sv"
`include "tmp/individual_1.sv"
`include "tmp/individual_2.sv"
`include "tmp/individual_3.sv"
`include "tmp/individual_4.sv"
`include "tmp/individual_5.sv"
`include "tmp/individual_6.sv"
`include "tmp/individual_7.sv"
`include "tmp/individual_8.sv"
`include "tmp/individual_9.sv"
`include "tmp/individual_10.sv"
`include "tmp/individual_11.sv"
`include "tmp/individual_12.sv"
`include "tmp/individual_13.sv"
`include "tmp/individual_14.sv"
`include "tmp/individual_15.sv"
`include "tmp/individual_16.sv"
`include "tmp/individual_17.sv"
`include "tmp/individual_18.sv"
`include "tmp/individual_19.sv"
`include "tmp/individual_20.sv"
`include "tmp/individual_21.sv"
`include "tmp/individual_22.sv"
`include "tmp/individual_23.sv"
`include "tmp/individual_24.sv"
`include "tmp/individual_25.sv"
`include "tmp/individual_26.sv"
`include "tmp/individual_27.sv"
`include "tmp/individual_28.sv"
`include "tmp/individual_29.sv"
`include "tmp/individual_30.sv"
`include "tmp/individual_31.sv"
`include "tmp/individual_32.sv"
`include "tmp/individual_33.sv"
`include "tmp/individual_34.sv"
`include "tmp/individual_35.sv"
`include "tmp/individual_36.sv"
`include "tmp/individual_37.sv"
`include "tmp/individual_38.sv"
`include "tmp/individual_39.sv"
`include "tmp/individual_40.sv"
`include "tmp/individual_41.sv"
`include "tmp/individual_42.sv"
`include "tmp/individual_43.sv"
`include "tmp/individual_44.sv"
`include "tmp/individual_45.sv"
`include "tmp/individual_46.sv"
`include "tmp/individual_47.sv"
`include "tmp/individual_48.sv"
`include "tmp/individual_49.sv"
`include "tmp/individual_50.sv"
`include "tmp/individual_51.sv"
`include "tmp/individual_52.sv"
`include "tmp/individual_53.sv"
`include "tmp/individual_54.sv"
`include "tmp/individual_55.sv"
`include "tmp/individual_56.sv"
`include "tmp/individual_57.sv"
`include "tmp/individual_58.sv"
`include "tmp/individual_59.sv"
`include "tmp/individual_60.sv"
`include "tmp/individual_61.sv"
`include "tmp/individual_62.sv"
`include "tmp/individual_63.sv"
`include "tmp/individual_64.sv"
`include "tmp/individual_65.sv"
`include "tmp/individual_66.sv"
`include "tmp/individual_67.sv"
`include "tmp/individual_68.sv"
`include "tmp/individual_69.sv"
`include "tmp/individual_70.sv"
`include "tmp/individual_71.sv"
`include "tmp/individual_72.sv"
`include "tmp/individual_73.sv"
`include "tmp/individual_74.sv"
`include "tmp/individual_75.sv"
`include "tmp/individual_76.sv"
`include "tmp/individual_77.sv"
`include "tmp/individual_78.sv"
`include "tmp/individual_79.sv"
`include "tmp/individual_80.sv"
`include "tmp/individual_81.sv"
`include "tmp/individual_82.sv"
`include "tmp/individual_83.sv"
`include "tmp/individual_84.sv"
`include "tmp/individual_85.sv"
`include "tmp/individual_86.sv"
`include "tmp/individual_87.sv"
`include "tmp/individual_88.sv"
`include "tmp/individual_89.sv"
`include "tmp/individual_90.sv"
`include "tmp/individual_91.sv"
`include "tmp/individual_92.sv"
`include "tmp/individual_93.sv"
`include "tmp/individual_94.sv"
`include "tmp/individual_95.sv"
`include "tmp/individual_96.sv"
`include "tmp/individual_97.sv"
`include "tmp/individual_98.sv"
`include "tmp/individual_99.sv"
`include "tmp/individual_100.sv"
`include "tmp/individual_101.sv"
`include "tmp/individual_102.sv"
`include "tmp/individual_103.sv"
`include "tmp/individual_104.sv"
`include "tmp/individual_105.sv"
`include "tmp/individual_106.sv"
`include "tmp/individual_107.sv"
`include "tmp/individual_108.sv"
`include "tmp/individual_109.sv"
`include "tmp/individual_110.sv"
`include "tmp/individual_111.sv"
`include "tmp/individual_112.sv"
`include "tmp/individual_113.sv"
`include "tmp/individual_114.sv"
`include "tmp/individual_115.sv"
`include "tmp/individual_116.sv"
`include "tmp/individual_117.sv"
`include "tmp/individual_118.sv"
`include "tmp/individual_119.sv"
`include "tmp/individual_120.sv"
`include "tmp/individual_121.sv"
`include "tmp/individual_122.sv"
`include "tmp/individual_123.sv"
`include "tmp/individual_124.sv"
`include "tmp/individual_125.sv"
`include "tmp/individual_126.sv"
`include "tmp/individual_127.sv"
`include "tmp/individual_128.sv"
`include "tmp/individual_129.sv"
`include "tmp/individual_130.sv"
`include "tmp/individual_131.sv"
`include "tmp/individual_132.sv"
`include "tmp/individual_133.sv"
`include "tmp/individual_134.sv"
`include "tmp/individual_135.sv"
`include "tmp/individual_136.sv"
`include "tmp/individual_137.sv"
`include "tmp/individual_138.sv"
`include "tmp/individual_139.sv"
`include "tmp/individual_140.sv"
`include "tmp/individual_141.sv"
`include "tmp/individual_142.sv"
`include "tmp/individual_143.sv"
`include "tmp/individual_144.sv"
`include "tmp/individual_145.sv"
`include "tmp/individual_146.sv"
`include "tmp/individual_147.sv"
`include "tmp/individual_148.sv"
`include "tmp/individual_149.sv"
`include "tmp/individual_150.sv"
`include "tmp/individual_151.sv"
`include "tmp/individual_152.sv"
`include "tmp/individual_153.sv"
`include "tmp/individual_154.sv"
`include "tmp/individual_155.sv"
`include "tmp/individual_156.sv"
`include "tmp/individual_157.sv"
`include "tmp/individual_158.sv"
`include "tmp/individual_159.sv"
`include "tmp/individual_160.sv"
`include "tmp/individual_161.sv"
`include "tmp/individual_162.sv"
`include "tmp/individual_163.sv"
`include "tmp/individual_164.sv"
`include "tmp/individual_165.sv"
`include "tmp/individual_166.sv"
`include "tmp/individual_167.sv"
`include "tmp/individual_168.sv"
`include "tmp/individual_169.sv"
`include "tmp/individual_170.sv"
`include "tmp/individual_171.sv"
`include "tmp/individual_172.sv"
`include "tmp/individual_173.sv"
`include "tmp/individual_174.sv"
`include "tmp/individual_175.sv"
`include "tmp/individual_176.sv"
`include "tmp/individual_177.sv"
`include "tmp/individual_178.sv"
`include "tmp/individual_179.sv"
`include "tmp/individual_180.sv"
`include "tmp/individual_181.sv"
`include "tmp/individual_182.sv"
`include "tmp/individual_183.sv"
`include "tmp/individual_184.sv"
`include "tmp/individual_185.sv"
`include "tmp/individual_186.sv"
`include "tmp/individual_187.sv"
`include "tmp/individual_188.sv"
`include "tmp/individual_189.sv"
`include "tmp/individual_190.sv"
`include "tmp/individual_191.sv"
`include "tmp/individual_192.sv"
`include "tmp/individual_193.sv"
`include "tmp/individual_194.sv"
`include "tmp/individual_195.sv"
`include "tmp/individual_196.sv"
`include "tmp/individual_197.sv"
`include "tmp/individual_198.sv"
`include "tmp/individual_199.sv"
`include "tmp/individual_200.sv"
`include "tmp/individual_201.sv"
`include "tmp/individual_202.sv"
`include "tmp/individual_203.sv"
`include "tmp/individual_204.sv"
`include "tmp/individual_205.sv"
`include "tmp/individual_206.sv"
`include "tmp/individual_207.sv"
`include "tmp/individual_208.sv"
`include "tmp/individual_209.sv"
`include "tmp/individual_210.sv"
`include "tmp/individual_211.sv"
`include "tmp/individual_212.sv"
`include "tmp/individual_213.sv"
`include "tmp/individual_214.sv"
`include "tmp/individual_215.sv"
`include "tmp/individual_216.sv"
`include "tmp/individual_217.sv"
`include "tmp/individual_218.sv"
`include "tmp/individual_219.sv"
`include "tmp/individual_220.sv"
`include "tmp/individual_221.sv"
`include "tmp/individual_222.sv"
`include "tmp/individual_223.sv"
`include "tmp/individual_224.sv"
`include "tmp/individual_225.sv"
`include "tmp/individual_226.sv"
`include "tmp/individual_227.sv"
`include "tmp/individual_228.sv"
`include "tmp/individual_229.sv"
`include "tmp/individual_230.sv"
`include "tmp/individual_231.sv"
`include "tmp/individual_232.sv"
`include "tmp/individual_233.sv"
`include "tmp/individual_234.sv"
`include "tmp/individual_235.sv"
`include "tmp/individual_236.sv"
`include "tmp/individual_237.sv"
`include "tmp/individual_238.sv"
`include "tmp/individual_239.sv"
`include "tmp/individual_240.sv"
`include "tmp/individual_241.sv"
`include "tmp/individual_242.sv"
`include "tmp/individual_243.sv"
`include "tmp/individual_244.sv"
`include "tmp/individual_245.sv"
`include "tmp/individual_246.sv"
`include "tmp/individual_247.sv"
`include "tmp/individual_248.sv"
`include "tmp/individual_249.sv"
`include "tmp/individual_250.sv"
`include "tmp/individual_251.sv"
`include "tmp/individual_252.sv"
`include "tmp/individual_253.sv"
`include "tmp/individual_254.sv"
`include "tmp/individual_255.sv"
`include "tmp/individual_256.sv"
`include "tmp/individual_257.sv"
`include "tmp/individual_258.sv"
`include "tmp/individual_259.sv"
`include "tmp/individual_260.sv"
`include "tmp/individual_261.sv"
`include "tmp/individual_262.sv"
`include "tmp/individual_263.sv"
`include "tmp/individual_264.sv"
`include "tmp/individual_265.sv"
`include "tmp/individual_266.sv"
`include "tmp/individual_267.sv"
`include "tmp/individual_268.sv"
`include "tmp/individual_269.sv"
`include "tmp/individual_270.sv"
`include "tmp/individual_271.sv"
`include "tmp/individual_272.sv"
`include "tmp/individual_273.sv"
`include "tmp/individual_274.sv"
`include "tmp/individual_275.sv"
`include "tmp/individual_276.sv"
`include "tmp/individual_277.sv"
`include "tmp/individual_278.sv"
`include "tmp/individual_279.sv"
`include "tmp/individual_280.sv"
`include "tmp/individual_281.sv"
`include "tmp/individual_282.sv"
`include "tmp/individual_283.sv"
`include "tmp/individual_284.sv"
`include "tmp/individual_285.sv"
`include "tmp/individual_286.sv"
`include "tmp/individual_287.sv"
`include "tmp/individual_288.sv"
`include "tmp/individual_289.sv"
`include "tmp/individual_290.sv"
`include "tmp/individual_291.sv"
`include "tmp/individual_292.sv"
`include "tmp/individual_293.sv"
`include "tmp/individual_294.sv"
`include "tmp/individual_295.sv"
`include "tmp/individual_296.sv"
`include "tmp/individual_297.sv"
`include "tmp/individual_298.sv"
`include "tmp/individual_299.sv"
`include "tmp/individual_300.sv"
`include "tmp/individual_301.sv"
`include "tmp/individual_302.sv"
`include "tmp/individual_303.sv"
`include "tmp/individual_304.sv"
`include "tmp/individual_305.sv"
`include "tmp/individual_306.sv"
`include "tmp/individual_307.sv"
`include "tmp/individual_308.sv"
`include "tmp/individual_309.sv"
`include "tmp/individual_310.sv"
`include "tmp/individual_311.sv"
`include "tmp/individual_312.sv"
`include "tmp/individual_313.sv"
`include "tmp/individual_314.sv"
`include "tmp/individual_315.sv"
`include "tmp/individual_316.sv"
`include "tmp/individual_317.sv"
`include "tmp/individual_318.sv"
`include "tmp/individual_319.sv"
`include "tmp/individual_320.sv"
`include "tmp/individual_321.sv"
`include "tmp/individual_322.sv"
`include "tmp/individual_323.sv"
`include "tmp/individual_324.sv"
`include "tmp/individual_325.sv"
`include "tmp/individual_326.sv"
`include "tmp/individual_327.sv"
`include "tmp/individual_328.sv"
`include "tmp/individual_329.sv"
`include "tmp/individual_330.sv"
`include "tmp/individual_331.sv"
`include "tmp/individual_332.sv"
`include "tmp/individual_333.sv"
`include "tmp/individual_334.sv"
`include "tmp/individual_335.sv"
`include "tmp/individual_336.sv"
`include "tmp/individual_337.sv"
`include "tmp/individual_338.sv"
`include "tmp/individual_339.sv"
`include "tmp/individual_340.sv"
`include "tmp/individual_341.sv"
`include "tmp/individual_342.sv"
`include "tmp/individual_343.sv"
`include "tmp/individual_344.sv"
`include "tmp/individual_345.sv"
`include "tmp/individual_346.sv"
`include "tmp/individual_347.sv"
`include "tmp/individual_348.sv"
`include "tmp/individual_349.sv"
`include "tmp/individual_350.sv"
`include "tmp/individual_351.sv"
`include "tmp/individual_352.sv"
`include "tmp/individual_353.sv"
`include "tmp/individual_354.sv"
`include "tmp/individual_355.sv"
`include "tmp/individual_356.sv"
`include "tmp/individual_357.sv"
`include "tmp/individual_358.sv"
`include "tmp/individual_359.sv"
`include "tmp/individual_360.sv"
`include "tmp/individual_361.sv"
`include "tmp/individual_362.sv"
`include "tmp/individual_363.sv"
`include "tmp/individual_364.sv"
`include "tmp/individual_365.sv"
`include "tmp/individual_366.sv"
`include "tmp/individual_367.sv"
`include "tmp/individual_368.sv"
`include "tmp/individual_369.sv"
`include "tmp/individual_370.sv"
`include "tmp/individual_371.sv"
`include "tmp/individual_372.sv"
`include "tmp/individual_373.sv"
`include "tmp/individual_374.sv"
`include "tmp/individual_375.sv"
`include "tmp/individual_376.sv"
`include "tmp/individual_377.sv"
`include "tmp/individual_378.sv"
`include "tmp/individual_379.sv"
`include "tmp/individual_380.sv"
`include "tmp/individual_381.sv"
`include "tmp/individual_382.sv"
`include "tmp/individual_383.sv"
`include "tmp/individual_384.sv"
`include "tmp/individual_385.sv"
`include "tmp/individual_386.sv"
`include "tmp/individual_387.sv"
`include "tmp/individual_388.sv"
`include "tmp/individual_389.sv"
`include "tmp/individual_390.sv"
`include "tmp/individual_391.sv"
`include "tmp/individual_392.sv"
`include "tmp/individual_393.sv"
`include "tmp/individual_394.sv"
`include "tmp/individual_395.sv"
`include "tmp/individual_396.sv"
`include "tmp/individual_397.sv"
`include "tmp/individual_398.sv"
`include "tmp/individual_399.sv"
`include "tmp/individual_400.sv"
`include "tmp/individual_401.sv"
`include "tmp/individual_402.sv"
`include "tmp/individual_403.sv"
`include "tmp/individual_404.sv"
`include "tmp/individual_405.sv"
`include "tmp/individual_406.sv"
`include "tmp/individual_407.sv"
`include "tmp/individual_408.sv"
`include "tmp/individual_409.sv"
`include "tmp/individual_410.sv"
`include "tmp/individual_411.sv"
`include "tmp/individual_412.sv"
`include "tmp/individual_413.sv"
`include "tmp/individual_414.sv"
`include "tmp/individual_415.sv"
`include "tmp/individual_416.sv"
`include "tmp/individual_417.sv"
`include "tmp/individual_418.sv"
`include "tmp/individual_419.sv"
`include "tmp/individual_420.sv"
`include "tmp/individual_421.sv"
`include "tmp/individual_422.sv"
`include "tmp/individual_423.sv"
`include "tmp/individual_424.sv"
`include "tmp/individual_425.sv"
`include "tmp/individual_426.sv"
`include "tmp/individual_427.sv"
`include "tmp/individual_428.sv"
`include "tmp/individual_429.sv"
`include "tmp/individual_430.sv"
`include "tmp/individual_431.sv"
`include "tmp/individual_432.sv"
`include "tmp/individual_433.sv"
`include "tmp/individual_434.sv"
`include "tmp/individual_435.sv"
`include "tmp/individual_436.sv"
`include "tmp/individual_437.sv"
`include "tmp/individual_438.sv"
`include "tmp/individual_439.sv"
`include "tmp/individual_440.sv"
`include "tmp/individual_441.sv"
`include "tmp/individual_442.sv"
`include "tmp/individual_443.sv"
`include "tmp/individual_444.sv"
`include "tmp/individual_445.sv"
`include "tmp/individual_446.sv"
`include "tmp/individual_447.sv"
`include "tmp/individual_448.sv"
`include "tmp/individual_449.sv"
`include "tmp/individual_450.sv"
`include "tmp/individual_451.sv"
`include "tmp/individual_452.sv"
`include "tmp/individual_453.sv"
`include "tmp/individual_454.sv"
`include "tmp/individual_455.sv"
`include "tmp/individual_456.sv"
`include "tmp/individual_457.sv"
`include "tmp/individual_458.sv"
`include "tmp/individual_459.sv"
`include "tmp/individual_460.sv"
`include "tmp/individual_461.sv"
`include "tmp/individual_462.sv"
`include "tmp/individual_463.sv"
`include "tmp/individual_464.sv"
`include "tmp/individual_465.sv"
`include "tmp/individual_466.sv"
`include "tmp/individual_467.sv"
`include "tmp/individual_468.sv"
`include "tmp/individual_469.sv"
`include "tmp/individual_470.sv"
`include "tmp/individual_471.sv"
`include "tmp/individual_472.sv"
`include "tmp/individual_473.sv"
`include "tmp/individual_474.sv"
`include "tmp/individual_475.sv"
`include "tmp/individual_476.sv"
`include "tmp/individual_477.sv"
`include "tmp/individual_478.sv"
`include "tmp/individual_479.sv"
`include "tmp/individual_480.sv"
`include "tmp/individual_481.sv"
`include "tmp/individual_482.sv"
`include "tmp/individual_483.sv"
`include "tmp/individual_484.sv"
`include "tmp/individual_485.sv"
`include "tmp/individual_486.sv"
`include "tmp/individual_487.sv"
`include "tmp/individual_488.sv"
`include "tmp/individual_489.sv"
`include "tmp/individual_490.sv"
`include "tmp/individual_491.sv"
`include "tmp/individual_492.sv"
`include "tmp/individual_493.sv"
`include "tmp/individual_494.sv"
`include "tmp/individual_495.sv"
`include "tmp/individual_496.sv"
`include "tmp/individual_497.sv"
`include "tmp/individual_498.sv"
`include "tmp/individual_499.sv"
`include "tmp/individual_500.sv"
`include "tmp/individual_501.sv"
`include "tmp/individual_502.sv"
`include "tmp/individual_503.sv"
`include "tmp/individual_504.sv"
`include "tmp/individual_505.sv"
`include "tmp/individual_506.sv"
`include "tmp/individual_507.sv"
`include "tmp/individual_508.sv"
`include "tmp/individual_509.sv"
`include "tmp/individual_510.sv"
`include "tmp/individual_511.sv"
`include "tmp/individual_512.sv"
`include "tmp/individual_513.sv"
`include "tmp/individual_514.sv"
`include "tmp/individual_515.sv"
`include "tmp/individual_516.sv"
`include "tmp/individual_517.sv"
`include "tmp/individual_518.sv"
`include "tmp/individual_519.sv"
`include "tmp/individual_520.sv"
`include "tmp/individual_521.sv"
`include "tmp/individual_522.sv"
`include "tmp/individual_523.sv"
`include "tmp/individual_524.sv"
`include "tmp/individual_525.sv"
`include "tmp/individual_526.sv"
`include "tmp/individual_527.sv"
`include "tmp/individual_528.sv"
`include "tmp/individual_529.sv"
`include "tmp/individual_530.sv"
`include "tmp/individual_531.sv"
`include "tmp/individual_532.sv"
`include "tmp/individual_533.sv"
`include "tmp/individual_534.sv"
`include "tmp/individual_535.sv"
`include "tmp/individual_536.sv"
`include "tmp/individual_537.sv"
`include "tmp/individual_538.sv"
`include "tmp/individual_539.sv"
`include "tmp/individual_540.sv"
`include "tmp/individual_541.sv"
`include "tmp/individual_542.sv"
`include "tmp/individual_543.sv"
`include "tmp/individual_544.sv"
`include "tmp/individual_545.sv"
`include "tmp/individual_546.sv"
`include "tmp/individual_547.sv"
`include "tmp/individual_548.sv"
`include "tmp/individual_549.sv"
`include "tmp/individual_550.sv"
`include "tmp/individual_551.sv"
`include "tmp/individual_552.sv"
`include "tmp/individual_553.sv"
`include "tmp/individual_554.sv"
`include "tmp/individual_555.sv"
`include "tmp/individual_556.sv"
`include "tmp/individual_557.sv"
`include "tmp/individual_558.sv"
`include "tmp/individual_559.sv"
`include "tmp/individual_560.sv"
`include "tmp/individual_561.sv"
`include "tmp/individual_562.sv"
`include "tmp/individual_563.sv"
`include "tmp/individual_564.sv"
`include "tmp/individual_565.sv"
`include "tmp/individual_566.sv"
`include "tmp/individual_567.sv"
`include "tmp/individual_568.sv"
`include "tmp/individual_569.sv"
`include "tmp/individual_570.sv"
`include "tmp/individual_571.sv"
`include "tmp/individual_572.sv"
`include "tmp/individual_573.sv"
`include "tmp/individual_574.sv"
`include "tmp/individual_575.sv"
`include "tmp/individual_576.sv"
`include "tmp/individual_577.sv"
`include "tmp/individual_578.sv"
`include "tmp/individual_579.sv"
`include "tmp/individual_580.sv"
`include "tmp/individual_581.sv"
`include "tmp/individual_582.sv"
`include "tmp/individual_583.sv"
`include "tmp/individual_584.sv"
`include "tmp/individual_585.sv"
`include "tmp/individual_586.sv"
`include "tmp/individual_587.sv"
`include "tmp/individual_588.sv"
`include "tmp/individual_589.sv"
`include "tmp/individual_590.sv"
`include "tmp/individual_591.sv"
`include "tmp/individual_592.sv"
`include "tmp/individual_593.sv"
`include "tmp/individual_594.sv"
`include "tmp/individual_595.sv"
`include "tmp/individual_596.sv"
`include "tmp/individual_597.sv"
`include "tmp/individual_598.sv"
`include "tmp/individual_599.sv"
`include "tmp/individual_600.sv"
`include "tmp/individual_601.sv"
`include "tmp/individual_602.sv"
`include "tmp/individual_603.sv"
`include "tmp/individual_604.sv"
`include "tmp/individual_605.sv"
`include "tmp/individual_606.sv"
`include "tmp/individual_607.sv"
`include "tmp/individual_608.sv"
`include "tmp/individual_609.sv"
`include "tmp/individual_610.sv"
`include "tmp/individual_611.sv"
`include "tmp/individual_612.sv"
`include "tmp/individual_613.sv"
`include "tmp/individual_614.sv"
`include "tmp/individual_615.sv"
`include "tmp/individual_616.sv"
`include "tmp/individual_617.sv"
`include "tmp/individual_618.sv"
`include "tmp/individual_619.sv"
`include "tmp/individual_620.sv"
`include "tmp/individual_621.sv"
`include "tmp/individual_622.sv"
`include "tmp/individual_623.sv"
`include "tmp/individual_624.sv"
`include "tmp/individual_625.sv"
`include "tmp/individual_626.sv"
`include "tmp/individual_627.sv"
`include "tmp/individual_628.sv"
`include "tmp/individual_629.sv"
`include "tmp/individual_630.sv"
`include "tmp/individual_631.sv"
`include "tmp/individual_632.sv"
`include "tmp/individual_633.sv"
`include "tmp/individual_634.sv"
`include "tmp/individual_635.sv"
`include "tmp/individual_636.sv"
`include "tmp/individual_637.sv"
`include "tmp/individual_638.sv"
`include "tmp/individual_639.sv"
`include "tmp/individual_640.sv"
`include "tmp/individual_641.sv"
`include "tmp/individual_642.sv"
`include "tmp/individual_643.sv"
`include "tmp/individual_644.sv"
`include "tmp/individual_645.sv"
`include "tmp/individual_646.sv"
`include "tmp/individual_647.sv"
`include "tmp/individual_648.sv"
`include "tmp/individual_649.sv"
`include "tmp/individual_650.sv"
`include "tmp/individual_651.sv"
`include "tmp/individual_652.sv"
`include "tmp/individual_653.sv"
`include "tmp/individual_654.sv"
`include "tmp/individual_655.sv"
`include "tmp/individual_656.sv"
`include "tmp/individual_657.sv"
`include "tmp/individual_658.sv"
`include "tmp/individual_659.sv"
`include "tmp/individual_660.sv"
`include "tmp/individual_661.sv"
`include "tmp/individual_662.sv"
`include "tmp/individual_663.sv"
`include "tmp/individual_664.sv"
`include "tmp/individual_665.sv"
`include "tmp/individual_666.sv"
`include "tmp/individual_667.sv"
`include "tmp/individual_668.sv"
`include "tmp/individual_669.sv"
`include "tmp/individual_670.sv"
`include "tmp/individual_671.sv"
`include "tmp/individual_672.sv"
`include "tmp/individual_673.sv"
`include "tmp/individual_674.sv"
`include "tmp/individual_675.sv"
`include "tmp/individual_676.sv"
`include "tmp/individual_677.sv"
`include "tmp/individual_678.sv"
`include "tmp/individual_679.sv"
`include "tmp/individual_680.sv"
`include "tmp/individual_681.sv"
`include "tmp/individual_682.sv"
`include "tmp/individual_683.sv"
`include "tmp/individual_684.sv"
`include "tmp/individual_685.sv"
`include "tmp/individual_686.sv"
`include "tmp/individual_687.sv"
`include "tmp/individual_688.sv"
`include "tmp/individual_689.sv"
`include "tmp/individual_690.sv"
`include "tmp/individual_691.sv"
`include "tmp/individual_692.sv"
`include "tmp/individual_693.sv"
`include "tmp/individual_694.sv"
`include "tmp/individual_695.sv"
`include "tmp/individual_696.sv"
`include "tmp/individual_697.sv"
`include "tmp/individual_698.sv"
`include "tmp/individual_699.sv"
`include "tmp/individual_700.sv"
`include "tmp/individual_701.sv"
`include "tmp/individual_702.sv"
`include "tmp/individual_703.sv"
`include "tmp/individual_704.sv"
`include "tmp/individual_705.sv"
`include "tmp/individual_706.sv"
`include "tmp/individual_707.sv"
`include "tmp/individual_708.sv"
`include "tmp/individual_709.sv"
`include "tmp/individual_710.sv"
`include "tmp/individual_711.sv"
`include "tmp/individual_712.sv"
`include "tmp/individual_713.sv"
`include "tmp/individual_714.sv"
`include "tmp/individual_715.sv"
`include "tmp/individual_716.sv"
`include "tmp/individual_717.sv"
`include "tmp/individual_718.sv"
`include "tmp/individual_719.sv"
`include "tmp/individual_720.sv"
`include "tmp/individual_721.sv"
`include "tmp/individual_722.sv"
`include "tmp/individual_723.sv"
`include "tmp/individual_724.sv"
`include "tmp/individual_725.sv"
`include "tmp/individual_726.sv"
`include "tmp/individual_727.sv"
`include "tmp/individual_728.sv"
`include "tmp/individual_729.sv"
`include "tmp/individual_730.sv"
`include "tmp/individual_731.sv"
`include "tmp/individual_732.sv"
`include "tmp/individual_733.sv"
`include "tmp/individual_734.sv"
`include "tmp/individual_735.sv"
`include "tmp/individual_736.sv"
`include "tmp/individual_737.sv"
`include "tmp/individual_738.sv"
`include "tmp/individual_739.sv"
`include "tmp/individual_740.sv"
`include "tmp/individual_741.sv"
`include "tmp/individual_742.sv"
`include "tmp/individual_743.sv"
`include "tmp/individual_744.sv"
`include "tmp/individual_745.sv"
`include "tmp/individual_746.sv"
`include "tmp/individual_747.sv"
`include "tmp/individual_748.sv"
`include "tmp/individual_749.sv"

// Definitions
`define POPULATION_SIZE 750
`define TEST_COUNT 2
`define PERIOD 10

// Use parameter to pass population size to testbench
module testbench();
  // Use integer array to store fitness for all individuals
  integer fitness[`POPULATION_SIZE];

  // Define inputs and outputs to connect to the individuals
  reg clk;
  reg rst;
  reg [15:0] y3_current[`POPULATION_SIZE];
  reg [15:0] y3_expected;
  reg [15:0] y2_current[`POPULATION_SIZE];
  reg [15:0] y2_expected;
  reg [15:0] y1_current[`POPULATION_SIZE];
  reg [15:0] y1_expected;
  reg [15:0] y0_current[`POPULATION_SIZE];
  reg [15:0] y0_expected;

	reg [15:0] a1;
	reg [15:0] a0;
	reg [15:0] b1;
	reg [15:0] b0;

	// Array of testvectors to store expected values
	reg [127:0] testvectors[0:(`TEST_COUNT-1)];
	integer vectornum = 0;

	// Instantiate all the individuals
  individual_0 dut_0(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[0]), .y2(y2_current[0]), .y1(y1_current[0]), .y0(y0_current[0]));
  individual_1 dut_1(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[1]), .y2(y2_current[1]), .y1(y1_current[1]), .y0(y0_current[1]));
  individual_2 dut_2(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[2]), .y2(y2_current[2]), .y1(y1_current[2]), .y0(y0_current[2]));
  individual_3 dut_3(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[3]), .y2(y2_current[3]), .y1(y1_current[3]), .y0(y0_current[3]));
  individual_4 dut_4(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[4]), .y2(y2_current[4]), .y1(y1_current[4]), .y0(y0_current[4]));
  individual_5 dut_5(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[5]), .y2(y2_current[5]), .y1(y1_current[5]), .y0(y0_current[5]));
  individual_6 dut_6(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[6]), .y2(y2_current[6]), .y1(y1_current[6]), .y0(y0_current[6]));
  individual_7 dut_7(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[7]), .y2(y2_current[7]), .y1(y1_current[7]), .y0(y0_current[7]));
  individual_8 dut_8(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[8]), .y2(y2_current[8]), .y1(y1_current[8]), .y0(y0_current[8]));
  individual_9 dut_9(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[9]), .y2(y2_current[9]), .y1(y1_current[9]), .y0(y0_current[9]));
  individual_10 dut_10(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[10]), .y2(y2_current[10]), .y1(y1_current[10]), .y0(y0_current[10]));
  individual_11 dut_11(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[11]), .y2(y2_current[11]), .y1(y1_current[11]), .y0(y0_current[11]));
  individual_12 dut_12(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[12]), .y2(y2_current[12]), .y1(y1_current[12]), .y0(y0_current[12]));
  individual_13 dut_13(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[13]), .y2(y2_current[13]), .y1(y1_current[13]), .y0(y0_current[13]));
  individual_14 dut_14(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[14]), .y2(y2_current[14]), .y1(y1_current[14]), .y0(y0_current[14]));
  individual_15 dut_15(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[15]), .y2(y2_current[15]), .y1(y1_current[15]), .y0(y0_current[15]));
  individual_16 dut_16(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[16]), .y2(y2_current[16]), .y1(y1_current[16]), .y0(y0_current[16]));
  individual_17 dut_17(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[17]), .y2(y2_current[17]), .y1(y1_current[17]), .y0(y0_current[17]));
  individual_18 dut_18(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[18]), .y2(y2_current[18]), .y1(y1_current[18]), .y0(y0_current[18]));
  individual_19 dut_19(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[19]), .y2(y2_current[19]), .y1(y1_current[19]), .y0(y0_current[19]));
  individual_20 dut_20(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[20]), .y2(y2_current[20]), .y1(y1_current[20]), .y0(y0_current[20]));
  individual_21 dut_21(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[21]), .y2(y2_current[21]), .y1(y1_current[21]), .y0(y0_current[21]));
  individual_22 dut_22(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[22]), .y2(y2_current[22]), .y1(y1_current[22]), .y0(y0_current[22]));
  individual_23 dut_23(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[23]), .y2(y2_current[23]), .y1(y1_current[23]), .y0(y0_current[23]));
  individual_24 dut_24(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[24]), .y2(y2_current[24]), .y1(y1_current[24]), .y0(y0_current[24]));
  individual_25 dut_25(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[25]), .y2(y2_current[25]), .y1(y1_current[25]), .y0(y0_current[25]));
  individual_26 dut_26(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[26]), .y2(y2_current[26]), .y1(y1_current[26]), .y0(y0_current[26]));
  individual_27 dut_27(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[27]), .y2(y2_current[27]), .y1(y1_current[27]), .y0(y0_current[27]));
  individual_28 dut_28(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[28]), .y2(y2_current[28]), .y1(y1_current[28]), .y0(y0_current[28]));
  individual_29 dut_29(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[29]), .y2(y2_current[29]), .y1(y1_current[29]), .y0(y0_current[29]));
  individual_30 dut_30(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[30]), .y2(y2_current[30]), .y1(y1_current[30]), .y0(y0_current[30]));
  individual_31 dut_31(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[31]), .y2(y2_current[31]), .y1(y1_current[31]), .y0(y0_current[31]));
  individual_32 dut_32(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[32]), .y2(y2_current[32]), .y1(y1_current[32]), .y0(y0_current[32]));
  individual_33 dut_33(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[33]), .y2(y2_current[33]), .y1(y1_current[33]), .y0(y0_current[33]));
  individual_34 dut_34(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[34]), .y2(y2_current[34]), .y1(y1_current[34]), .y0(y0_current[34]));
  individual_35 dut_35(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[35]), .y2(y2_current[35]), .y1(y1_current[35]), .y0(y0_current[35]));
  individual_36 dut_36(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[36]), .y2(y2_current[36]), .y1(y1_current[36]), .y0(y0_current[36]));
  individual_37 dut_37(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[37]), .y2(y2_current[37]), .y1(y1_current[37]), .y0(y0_current[37]));
  individual_38 dut_38(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[38]), .y2(y2_current[38]), .y1(y1_current[38]), .y0(y0_current[38]));
  individual_39 dut_39(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[39]), .y2(y2_current[39]), .y1(y1_current[39]), .y0(y0_current[39]));
  individual_40 dut_40(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[40]), .y2(y2_current[40]), .y1(y1_current[40]), .y0(y0_current[40]));
  individual_41 dut_41(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[41]), .y2(y2_current[41]), .y1(y1_current[41]), .y0(y0_current[41]));
  individual_42 dut_42(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[42]), .y2(y2_current[42]), .y1(y1_current[42]), .y0(y0_current[42]));
  individual_43 dut_43(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[43]), .y2(y2_current[43]), .y1(y1_current[43]), .y0(y0_current[43]));
  individual_44 dut_44(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[44]), .y2(y2_current[44]), .y1(y1_current[44]), .y0(y0_current[44]));
  individual_45 dut_45(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[45]), .y2(y2_current[45]), .y1(y1_current[45]), .y0(y0_current[45]));
  individual_46 dut_46(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[46]), .y2(y2_current[46]), .y1(y1_current[46]), .y0(y0_current[46]));
  individual_47 dut_47(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[47]), .y2(y2_current[47]), .y1(y1_current[47]), .y0(y0_current[47]));
  individual_48 dut_48(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[48]), .y2(y2_current[48]), .y1(y1_current[48]), .y0(y0_current[48]));
  individual_49 dut_49(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[49]), .y2(y2_current[49]), .y1(y1_current[49]), .y0(y0_current[49]));
  individual_50 dut_50(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[50]), .y2(y2_current[50]), .y1(y1_current[50]), .y0(y0_current[50]));
  individual_51 dut_51(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[51]), .y2(y2_current[51]), .y1(y1_current[51]), .y0(y0_current[51]));
  individual_52 dut_52(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[52]), .y2(y2_current[52]), .y1(y1_current[52]), .y0(y0_current[52]));
  individual_53 dut_53(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[53]), .y2(y2_current[53]), .y1(y1_current[53]), .y0(y0_current[53]));
  individual_54 dut_54(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[54]), .y2(y2_current[54]), .y1(y1_current[54]), .y0(y0_current[54]));
  individual_55 dut_55(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[55]), .y2(y2_current[55]), .y1(y1_current[55]), .y0(y0_current[55]));
  individual_56 dut_56(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[56]), .y2(y2_current[56]), .y1(y1_current[56]), .y0(y0_current[56]));
  individual_57 dut_57(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[57]), .y2(y2_current[57]), .y1(y1_current[57]), .y0(y0_current[57]));
  individual_58 dut_58(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[58]), .y2(y2_current[58]), .y1(y1_current[58]), .y0(y0_current[58]));
  individual_59 dut_59(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[59]), .y2(y2_current[59]), .y1(y1_current[59]), .y0(y0_current[59]));
  individual_60 dut_60(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[60]), .y2(y2_current[60]), .y1(y1_current[60]), .y0(y0_current[60]));
  individual_61 dut_61(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[61]), .y2(y2_current[61]), .y1(y1_current[61]), .y0(y0_current[61]));
  individual_62 dut_62(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[62]), .y2(y2_current[62]), .y1(y1_current[62]), .y0(y0_current[62]));
  individual_63 dut_63(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[63]), .y2(y2_current[63]), .y1(y1_current[63]), .y0(y0_current[63]));
  individual_64 dut_64(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[64]), .y2(y2_current[64]), .y1(y1_current[64]), .y0(y0_current[64]));
  individual_65 dut_65(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[65]), .y2(y2_current[65]), .y1(y1_current[65]), .y0(y0_current[65]));
  individual_66 dut_66(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[66]), .y2(y2_current[66]), .y1(y1_current[66]), .y0(y0_current[66]));
  individual_67 dut_67(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[67]), .y2(y2_current[67]), .y1(y1_current[67]), .y0(y0_current[67]));
  individual_68 dut_68(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[68]), .y2(y2_current[68]), .y1(y1_current[68]), .y0(y0_current[68]));
  individual_69 dut_69(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[69]), .y2(y2_current[69]), .y1(y1_current[69]), .y0(y0_current[69]));
  individual_70 dut_70(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[70]), .y2(y2_current[70]), .y1(y1_current[70]), .y0(y0_current[70]));
  individual_71 dut_71(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[71]), .y2(y2_current[71]), .y1(y1_current[71]), .y0(y0_current[71]));
  individual_72 dut_72(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[72]), .y2(y2_current[72]), .y1(y1_current[72]), .y0(y0_current[72]));
  individual_73 dut_73(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[73]), .y2(y2_current[73]), .y1(y1_current[73]), .y0(y0_current[73]));
  individual_74 dut_74(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[74]), .y2(y2_current[74]), .y1(y1_current[74]), .y0(y0_current[74]));
  individual_75 dut_75(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[75]), .y2(y2_current[75]), .y1(y1_current[75]), .y0(y0_current[75]));
  individual_76 dut_76(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[76]), .y2(y2_current[76]), .y1(y1_current[76]), .y0(y0_current[76]));
  individual_77 dut_77(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[77]), .y2(y2_current[77]), .y1(y1_current[77]), .y0(y0_current[77]));
  individual_78 dut_78(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[78]), .y2(y2_current[78]), .y1(y1_current[78]), .y0(y0_current[78]));
  individual_79 dut_79(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[79]), .y2(y2_current[79]), .y1(y1_current[79]), .y0(y0_current[79]));
  individual_80 dut_80(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[80]), .y2(y2_current[80]), .y1(y1_current[80]), .y0(y0_current[80]));
  individual_81 dut_81(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[81]), .y2(y2_current[81]), .y1(y1_current[81]), .y0(y0_current[81]));
  individual_82 dut_82(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[82]), .y2(y2_current[82]), .y1(y1_current[82]), .y0(y0_current[82]));
  individual_83 dut_83(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[83]), .y2(y2_current[83]), .y1(y1_current[83]), .y0(y0_current[83]));
  individual_84 dut_84(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[84]), .y2(y2_current[84]), .y1(y1_current[84]), .y0(y0_current[84]));
  individual_85 dut_85(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[85]), .y2(y2_current[85]), .y1(y1_current[85]), .y0(y0_current[85]));
  individual_86 dut_86(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[86]), .y2(y2_current[86]), .y1(y1_current[86]), .y0(y0_current[86]));
  individual_87 dut_87(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[87]), .y2(y2_current[87]), .y1(y1_current[87]), .y0(y0_current[87]));
  individual_88 dut_88(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[88]), .y2(y2_current[88]), .y1(y1_current[88]), .y0(y0_current[88]));
  individual_89 dut_89(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[89]), .y2(y2_current[89]), .y1(y1_current[89]), .y0(y0_current[89]));
  individual_90 dut_90(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[90]), .y2(y2_current[90]), .y1(y1_current[90]), .y0(y0_current[90]));
  individual_91 dut_91(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[91]), .y2(y2_current[91]), .y1(y1_current[91]), .y0(y0_current[91]));
  individual_92 dut_92(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[92]), .y2(y2_current[92]), .y1(y1_current[92]), .y0(y0_current[92]));
  individual_93 dut_93(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[93]), .y2(y2_current[93]), .y1(y1_current[93]), .y0(y0_current[93]));
  individual_94 dut_94(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[94]), .y2(y2_current[94]), .y1(y1_current[94]), .y0(y0_current[94]));
  individual_95 dut_95(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[95]), .y2(y2_current[95]), .y1(y1_current[95]), .y0(y0_current[95]));
  individual_96 dut_96(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[96]), .y2(y2_current[96]), .y1(y1_current[96]), .y0(y0_current[96]));
  individual_97 dut_97(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[97]), .y2(y2_current[97]), .y1(y1_current[97]), .y0(y0_current[97]));
  individual_98 dut_98(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[98]), .y2(y2_current[98]), .y1(y1_current[98]), .y0(y0_current[98]));
  individual_99 dut_99(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[99]), .y2(y2_current[99]), .y1(y1_current[99]), .y0(y0_current[99]));
  individual_100 dut_100(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[100]), .y2(y2_current[100]), .y1(y1_current[100]), .y0(y0_current[100]));
  individual_101 dut_101(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[101]), .y2(y2_current[101]), .y1(y1_current[101]), .y0(y0_current[101]));
  individual_102 dut_102(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[102]), .y2(y2_current[102]), .y1(y1_current[102]), .y0(y0_current[102]));
  individual_103 dut_103(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[103]), .y2(y2_current[103]), .y1(y1_current[103]), .y0(y0_current[103]));
  individual_104 dut_104(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[104]), .y2(y2_current[104]), .y1(y1_current[104]), .y0(y0_current[104]));
  individual_105 dut_105(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[105]), .y2(y2_current[105]), .y1(y1_current[105]), .y0(y0_current[105]));
  individual_106 dut_106(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[106]), .y2(y2_current[106]), .y1(y1_current[106]), .y0(y0_current[106]));
  individual_107 dut_107(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[107]), .y2(y2_current[107]), .y1(y1_current[107]), .y0(y0_current[107]));
  individual_108 dut_108(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[108]), .y2(y2_current[108]), .y1(y1_current[108]), .y0(y0_current[108]));
  individual_109 dut_109(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[109]), .y2(y2_current[109]), .y1(y1_current[109]), .y0(y0_current[109]));
  individual_110 dut_110(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[110]), .y2(y2_current[110]), .y1(y1_current[110]), .y0(y0_current[110]));
  individual_111 dut_111(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[111]), .y2(y2_current[111]), .y1(y1_current[111]), .y0(y0_current[111]));
  individual_112 dut_112(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[112]), .y2(y2_current[112]), .y1(y1_current[112]), .y0(y0_current[112]));
  individual_113 dut_113(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[113]), .y2(y2_current[113]), .y1(y1_current[113]), .y0(y0_current[113]));
  individual_114 dut_114(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[114]), .y2(y2_current[114]), .y1(y1_current[114]), .y0(y0_current[114]));
  individual_115 dut_115(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[115]), .y2(y2_current[115]), .y1(y1_current[115]), .y0(y0_current[115]));
  individual_116 dut_116(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[116]), .y2(y2_current[116]), .y1(y1_current[116]), .y0(y0_current[116]));
  individual_117 dut_117(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[117]), .y2(y2_current[117]), .y1(y1_current[117]), .y0(y0_current[117]));
  individual_118 dut_118(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[118]), .y2(y2_current[118]), .y1(y1_current[118]), .y0(y0_current[118]));
  individual_119 dut_119(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[119]), .y2(y2_current[119]), .y1(y1_current[119]), .y0(y0_current[119]));
  individual_120 dut_120(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[120]), .y2(y2_current[120]), .y1(y1_current[120]), .y0(y0_current[120]));
  individual_121 dut_121(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[121]), .y2(y2_current[121]), .y1(y1_current[121]), .y0(y0_current[121]));
  individual_122 dut_122(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[122]), .y2(y2_current[122]), .y1(y1_current[122]), .y0(y0_current[122]));
  individual_123 dut_123(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[123]), .y2(y2_current[123]), .y1(y1_current[123]), .y0(y0_current[123]));
  individual_124 dut_124(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[124]), .y2(y2_current[124]), .y1(y1_current[124]), .y0(y0_current[124]));
  individual_125 dut_125(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[125]), .y2(y2_current[125]), .y1(y1_current[125]), .y0(y0_current[125]));
  individual_126 dut_126(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[126]), .y2(y2_current[126]), .y1(y1_current[126]), .y0(y0_current[126]));
  individual_127 dut_127(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[127]), .y2(y2_current[127]), .y1(y1_current[127]), .y0(y0_current[127]));
  individual_128 dut_128(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[128]), .y2(y2_current[128]), .y1(y1_current[128]), .y0(y0_current[128]));
  individual_129 dut_129(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[129]), .y2(y2_current[129]), .y1(y1_current[129]), .y0(y0_current[129]));
  individual_130 dut_130(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[130]), .y2(y2_current[130]), .y1(y1_current[130]), .y0(y0_current[130]));
  individual_131 dut_131(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[131]), .y2(y2_current[131]), .y1(y1_current[131]), .y0(y0_current[131]));
  individual_132 dut_132(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[132]), .y2(y2_current[132]), .y1(y1_current[132]), .y0(y0_current[132]));
  individual_133 dut_133(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[133]), .y2(y2_current[133]), .y1(y1_current[133]), .y0(y0_current[133]));
  individual_134 dut_134(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[134]), .y2(y2_current[134]), .y1(y1_current[134]), .y0(y0_current[134]));
  individual_135 dut_135(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[135]), .y2(y2_current[135]), .y1(y1_current[135]), .y0(y0_current[135]));
  individual_136 dut_136(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[136]), .y2(y2_current[136]), .y1(y1_current[136]), .y0(y0_current[136]));
  individual_137 dut_137(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[137]), .y2(y2_current[137]), .y1(y1_current[137]), .y0(y0_current[137]));
  individual_138 dut_138(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[138]), .y2(y2_current[138]), .y1(y1_current[138]), .y0(y0_current[138]));
  individual_139 dut_139(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[139]), .y2(y2_current[139]), .y1(y1_current[139]), .y0(y0_current[139]));
  individual_140 dut_140(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[140]), .y2(y2_current[140]), .y1(y1_current[140]), .y0(y0_current[140]));
  individual_141 dut_141(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[141]), .y2(y2_current[141]), .y1(y1_current[141]), .y0(y0_current[141]));
  individual_142 dut_142(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[142]), .y2(y2_current[142]), .y1(y1_current[142]), .y0(y0_current[142]));
  individual_143 dut_143(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[143]), .y2(y2_current[143]), .y1(y1_current[143]), .y0(y0_current[143]));
  individual_144 dut_144(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[144]), .y2(y2_current[144]), .y1(y1_current[144]), .y0(y0_current[144]));
  individual_145 dut_145(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[145]), .y2(y2_current[145]), .y1(y1_current[145]), .y0(y0_current[145]));
  individual_146 dut_146(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[146]), .y2(y2_current[146]), .y1(y1_current[146]), .y0(y0_current[146]));
  individual_147 dut_147(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[147]), .y2(y2_current[147]), .y1(y1_current[147]), .y0(y0_current[147]));
  individual_148 dut_148(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[148]), .y2(y2_current[148]), .y1(y1_current[148]), .y0(y0_current[148]));
  individual_149 dut_149(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[149]), .y2(y2_current[149]), .y1(y1_current[149]), .y0(y0_current[149]));
  individual_150 dut_150(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[150]), .y2(y2_current[150]), .y1(y1_current[150]), .y0(y0_current[150]));
  individual_151 dut_151(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[151]), .y2(y2_current[151]), .y1(y1_current[151]), .y0(y0_current[151]));
  individual_152 dut_152(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[152]), .y2(y2_current[152]), .y1(y1_current[152]), .y0(y0_current[152]));
  individual_153 dut_153(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[153]), .y2(y2_current[153]), .y1(y1_current[153]), .y0(y0_current[153]));
  individual_154 dut_154(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[154]), .y2(y2_current[154]), .y1(y1_current[154]), .y0(y0_current[154]));
  individual_155 dut_155(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[155]), .y2(y2_current[155]), .y1(y1_current[155]), .y0(y0_current[155]));
  individual_156 dut_156(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[156]), .y2(y2_current[156]), .y1(y1_current[156]), .y0(y0_current[156]));
  individual_157 dut_157(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[157]), .y2(y2_current[157]), .y1(y1_current[157]), .y0(y0_current[157]));
  individual_158 dut_158(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[158]), .y2(y2_current[158]), .y1(y1_current[158]), .y0(y0_current[158]));
  individual_159 dut_159(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[159]), .y2(y2_current[159]), .y1(y1_current[159]), .y0(y0_current[159]));
  individual_160 dut_160(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[160]), .y2(y2_current[160]), .y1(y1_current[160]), .y0(y0_current[160]));
  individual_161 dut_161(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[161]), .y2(y2_current[161]), .y1(y1_current[161]), .y0(y0_current[161]));
  individual_162 dut_162(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[162]), .y2(y2_current[162]), .y1(y1_current[162]), .y0(y0_current[162]));
  individual_163 dut_163(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[163]), .y2(y2_current[163]), .y1(y1_current[163]), .y0(y0_current[163]));
  individual_164 dut_164(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[164]), .y2(y2_current[164]), .y1(y1_current[164]), .y0(y0_current[164]));
  individual_165 dut_165(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[165]), .y2(y2_current[165]), .y1(y1_current[165]), .y0(y0_current[165]));
  individual_166 dut_166(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[166]), .y2(y2_current[166]), .y1(y1_current[166]), .y0(y0_current[166]));
  individual_167 dut_167(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[167]), .y2(y2_current[167]), .y1(y1_current[167]), .y0(y0_current[167]));
  individual_168 dut_168(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[168]), .y2(y2_current[168]), .y1(y1_current[168]), .y0(y0_current[168]));
  individual_169 dut_169(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[169]), .y2(y2_current[169]), .y1(y1_current[169]), .y0(y0_current[169]));
  individual_170 dut_170(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[170]), .y2(y2_current[170]), .y1(y1_current[170]), .y0(y0_current[170]));
  individual_171 dut_171(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[171]), .y2(y2_current[171]), .y1(y1_current[171]), .y0(y0_current[171]));
  individual_172 dut_172(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[172]), .y2(y2_current[172]), .y1(y1_current[172]), .y0(y0_current[172]));
  individual_173 dut_173(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[173]), .y2(y2_current[173]), .y1(y1_current[173]), .y0(y0_current[173]));
  individual_174 dut_174(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[174]), .y2(y2_current[174]), .y1(y1_current[174]), .y0(y0_current[174]));
  individual_175 dut_175(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[175]), .y2(y2_current[175]), .y1(y1_current[175]), .y0(y0_current[175]));
  individual_176 dut_176(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[176]), .y2(y2_current[176]), .y1(y1_current[176]), .y0(y0_current[176]));
  individual_177 dut_177(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[177]), .y2(y2_current[177]), .y1(y1_current[177]), .y0(y0_current[177]));
  individual_178 dut_178(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[178]), .y2(y2_current[178]), .y1(y1_current[178]), .y0(y0_current[178]));
  individual_179 dut_179(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[179]), .y2(y2_current[179]), .y1(y1_current[179]), .y0(y0_current[179]));
  individual_180 dut_180(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[180]), .y2(y2_current[180]), .y1(y1_current[180]), .y0(y0_current[180]));
  individual_181 dut_181(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[181]), .y2(y2_current[181]), .y1(y1_current[181]), .y0(y0_current[181]));
  individual_182 dut_182(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[182]), .y2(y2_current[182]), .y1(y1_current[182]), .y0(y0_current[182]));
  individual_183 dut_183(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[183]), .y2(y2_current[183]), .y1(y1_current[183]), .y0(y0_current[183]));
  individual_184 dut_184(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[184]), .y2(y2_current[184]), .y1(y1_current[184]), .y0(y0_current[184]));
  individual_185 dut_185(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[185]), .y2(y2_current[185]), .y1(y1_current[185]), .y0(y0_current[185]));
  individual_186 dut_186(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[186]), .y2(y2_current[186]), .y1(y1_current[186]), .y0(y0_current[186]));
  individual_187 dut_187(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[187]), .y2(y2_current[187]), .y1(y1_current[187]), .y0(y0_current[187]));
  individual_188 dut_188(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[188]), .y2(y2_current[188]), .y1(y1_current[188]), .y0(y0_current[188]));
  individual_189 dut_189(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[189]), .y2(y2_current[189]), .y1(y1_current[189]), .y0(y0_current[189]));
  individual_190 dut_190(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[190]), .y2(y2_current[190]), .y1(y1_current[190]), .y0(y0_current[190]));
  individual_191 dut_191(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[191]), .y2(y2_current[191]), .y1(y1_current[191]), .y0(y0_current[191]));
  individual_192 dut_192(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[192]), .y2(y2_current[192]), .y1(y1_current[192]), .y0(y0_current[192]));
  individual_193 dut_193(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[193]), .y2(y2_current[193]), .y1(y1_current[193]), .y0(y0_current[193]));
  individual_194 dut_194(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[194]), .y2(y2_current[194]), .y1(y1_current[194]), .y0(y0_current[194]));
  individual_195 dut_195(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[195]), .y2(y2_current[195]), .y1(y1_current[195]), .y0(y0_current[195]));
  individual_196 dut_196(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[196]), .y2(y2_current[196]), .y1(y1_current[196]), .y0(y0_current[196]));
  individual_197 dut_197(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[197]), .y2(y2_current[197]), .y1(y1_current[197]), .y0(y0_current[197]));
  individual_198 dut_198(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[198]), .y2(y2_current[198]), .y1(y1_current[198]), .y0(y0_current[198]));
  individual_199 dut_199(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[199]), .y2(y2_current[199]), .y1(y1_current[199]), .y0(y0_current[199]));
  individual_200 dut_200(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[200]), .y2(y2_current[200]), .y1(y1_current[200]), .y0(y0_current[200]));
  individual_201 dut_201(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[201]), .y2(y2_current[201]), .y1(y1_current[201]), .y0(y0_current[201]));
  individual_202 dut_202(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[202]), .y2(y2_current[202]), .y1(y1_current[202]), .y0(y0_current[202]));
  individual_203 dut_203(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[203]), .y2(y2_current[203]), .y1(y1_current[203]), .y0(y0_current[203]));
  individual_204 dut_204(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[204]), .y2(y2_current[204]), .y1(y1_current[204]), .y0(y0_current[204]));
  individual_205 dut_205(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[205]), .y2(y2_current[205]), .y1(y1_current[205]), .y0(y0_current[205]));
  individual_206 dut_206(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[206]), .y2(y2_current[206]), .y1(y1_current[206]), .y0(y0_current[206]));
  individual_207 dut_207(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[207]), .y2(y2_current[207]), .y1(y1_current[207]), .y0(y0_current[207]));
  individual_208 dut_208(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[208]), .y2(y2_current[208]), .y1(y1_current[208]), .y0(y0_current[208]));
  individual_209 dut_209(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[209]), .y2(y2_current[209]), .y1(y1_current[209]), .y0(y0_current[209]));
  individual_210 dut_210(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[210]), .y2(y2_current[210]), .y1(y1_current[210]), .y0(y0_current[210]));
  individual_211 dut_211(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[211]), .y2(y2_current[211]), .y1(y1_current[211]), .y0(y0_current[211]));
  individual_212 dut_212(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[212]), .y2(y2_current[212]), .y1(y1_current[212]), .y0(y0_current[212]));
  individual_213 dut_213(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[213]), .y2(y2_current[213]), .y1(y1_current[213]), .y0(y0_current[213]));
  individual_214 dut_214(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[214]), .y2(y2_current[214]), .y1(y1_current[214]), .y0(y0_current[214]));
  individual_215 dut_215(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[215]), .y2(y2_current[215]), .y1(y1_current[215]), .y0(y0_current[215]));
  individual_216 dut_216(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[216]), .y2(y2_current[216]), .y1(y1_current[216]), .y0(y0_current[216]));
  individual_217 dut_217(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[217]), .y2(y2_current[217]), .y1(y1_current[217]), .y0(y0_current[217]));
  individual_218 dut_218(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[218]), .y2(y2_current[218]), .y1(y1_current[218]), .y0(y0_current[218]));
  individual_219 dut_219(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[219]), .y2(y2_current[219]), .y1(y1_current[219]), .y0(y0_current[219]));
  individual_220 dut_220(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[220]), .y2(y2_current[220]), .y1(y1_current[220]), .y0(y0_current[220]));
  individual_221 dut_221(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[221]), .y2(y2_current[221]), .y1(y1_current[221]), .y0(y0_current[221]));
  individual_222 dut_222(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[222]), .y2(y2_current[222]), .y1(y1_current[222]), .y0(y0_current[222]));
  individual_223 dut_223(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[223]), .y2(y2_current[223]), .y1(y1_current[223]), .y0(y0_current[223]));
  individual_224 dut_224(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[224]), .y2(y2_current[224]), .y1(y1_current[224]), .y0(y0_current[224]));
  individual_225 dut_225(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[225]), .y2(y2_current[225]), .y1(y1_current[225]), .y0(y0_current[225]));
  individual_226 dut_226(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[226]), .y2(y2_current[226]), .y1(y1_current[226]), .y0(y0_current[226]));
  individual_227 dut_227(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[227]), .y2(y2_current[227]), .y1(y1_current[227]), .y0(y0_current[227]));
  individual_228 dut_228(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[228]), .y2(y2_current[228]), .y1(y1_current[228]), .y0(y0_current[228]));
  individual_229 dut_229(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[229]), .y2(y2_current[229]), .y1(y1_current[229]), .y0(y0_current[229]));
  individual_230 dut_230(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[230]), .y2(y2_current[230]), .y1(y1_current[230]), .y0(y0_current[230]));
  individual_231 dut_231(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[231]), .y2(y2_current[231]), .y1(y1_current[231]), .y0(y0_current[231]));
  individual_232 dut_232(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[232]), .y2(y2_current[232]), .y1(y1_current[232]), .y0(y0_current[232]));
  individual_233 dut_233(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[233]), .y2(y2_current[233]), .y1(y1_current[233]), .y0(y0_current[233]));
  individual_234 dut_234(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[234]), .y2(y2_current[234]), .y1(y1_current[234]), .y0(y0_current[234]));
  individual_235 dut_235(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[235]), .y2(y2_current[235]), .y1(y1_current[235]), .y0(y0_current[235]));
  individual_236 dut_236(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[236]), .y2(y2_current[236]), .y1(y1_current[236]), .y0(y0_current[236]));
  individual_237 dut_237(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[237]), .y2(y2_current[237]), .y1(y1_current[237]), .y0(y0_current[237]));
  individual_238 dut_238(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[238]), .y2(y2_current[238]), .y1(y1_current[238]), .y0(y0_current[238]));
  individual_239 dut_239(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[239]), .y2(y2_current[239]), .y1(y1_current[239]), .y0(y0_current[239]));
  individual_240 dut_240(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[240]), .y2(y2_current[240]), .y1(y1_current[240]), .y0(y0_current[240]));
  individual_241 dut_241(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[241]), .y2(y2_current[241]), .y1(y1_current[241]), .y0(y0_current[241]));
  individual_242 dut_242(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[242]), .y2(y2_current[242]), .y1(y1_current[242]), .y0(y0_current[242]));
  individual_243 dut_243(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[243]), .y2(y2_current[243]), .y1(y1_current[243]), .y0(y0_current[243]));
  individual_244 dut_244(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[244]), .y2(y2_current[244]), .y1(y1_current[244]), .y0(y0_current[244]));
  individual_245 dut_245(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[245]), .y2(y2_current[245]), .y1(y1_current[245]), .y0(y0_current[245]));
  individual_246 dut_246(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[246]), .y2(y2_current[246]), .y1(y1_current[246]), .y0(y0_current[246]));
  individual_247 dut_247(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[247]), .y2(y2_current[247]), .y1(y1_current[247]), .y0(y0_current[247]));
  individual_248 dut_248(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[248]), .y2(y2_current[248]), .y1(y1_current[248]), .y0(y0_current[248]));
  individual_249 dut_249(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[249]), .y2(y2_current[249]), .y1(y1_current[249]), .y0(y0_current[249]));
  individual_250 dut_250(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[250]), .y2(y2_current[250]), .y1(y1_current[250]), .y0(y0_current[250]));
  individual_251 dut_251(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[251]), .y2(y2_current[251]), .y1(y1_current[251]), .y0(y0_current[251]));
  individual_252 dut_252(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[252]), .y2(y2_current[252]), .y1(y1_current[252]), .y0(y0_current[252]));
  individual_253 dut_253(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[253]), .y2(y2_current[253]), .y1(y1_current[253]), .y0(y0_current[253]));
  individual_254 dut_254(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[254]), .y2(y2_current[254]), .y1(y1_current[254]), .y0(y0_current[254]));
  individual_255 dut_255(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[255]), .y2(y2_current[255]), .y1(y1_current[255]), .y0(y0_current[255]));
  individual_256 dut_256(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[256]), .y2(y2_current[256]), .y1(y1_current[256]), .y0(y0_current[256]));
  individual_257 dut_257(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[257]), .y2(y2_current[257]), .y1(y1_current[257]), .y0(y0_current[257]));
  individual_258 dut_258(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[258]), .y2(y2_current[258]), .y1(y1_current[258]), .y0(y0_current[258]));
  individual_259 dut_259(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[259]), .y2(y2_current[259]), .y1(y1_current[259]), .y0(y0_current[259]));
  individual_260 dut_260(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[260]), .y2(y2_current[260]), .y1(y1_current[260]), .y0(y0_current[260]));
  individual_261 dut_261(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[261]), .y2(y2_current[261]), .y1(y1_current[261]), .y0(y0_current[261]));
  individual_262 dut_262(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[262]), .y2(y2_current[262]), .y1(y1_current[262]), .y0(y0_current[262]));
  individual_263 dut_263(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[263]), .y2(y2_current[263]), .y1(y1_current[263]), .y0(y0_current[263]));
  individual_264 dut_264(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[264]), .y2(y2_current[264]), .y1(y1_current[264]), .y0(y0_current[264]));
  individual_265 dut_265(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[265]), .y2(y2_current[265]), .y1(y1_current[265]), .y0(y0_current[265]));
  individual_266 dut_266(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[266]), .y2(y2_current[266]), .y1(y1_current[266]), .y0(y0_current[266]));
  individual_267 dut_267(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[267]), .y2(y2_current[267]), .y1(y1_current[267]), .y0(y0_current[267]));
  individual_268 dut_268(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[268]), .y2(y2_current[268]), .y1(y1_current[268]), .y0(y0_current[268]));
  individual_269 dut_269(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[269]), .y2(y2_current[269]), .y1(y1_current[269]), .y0(y0_current[269]));
  individual_270 dut_270(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[270]), .y2(y2_current[270]), .y1(y1_current[270]), .y0(y0_current[270]));
  individual_271 dut_271(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[271]), .y2(y2_current[271]), .y1(y1_current[271]), .y0(y0_current[271]));
  individual_272 dut_272(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[272]), .y2(y2_current[272]), .y1(y1_current[272]), .y0(y0_current[272]));
  individual_273 dut_273(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[273]), .y2(y2_current[273]), .y1(y1_current[273]), .y0(y0_current[273]));
  individual_274 dut_274(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[274]), .y2(y2_current[274]), .y1(y1_current[274]), .y0(y0_current[274]));
  individual_275 dut_275(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[275]), .y2(y2_current[275]), .y1(y1_current[275]), .y0(y0_current[275]));
  individual_276 dut_276(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[276]), .y2(y2_current[276]), .y1(y1_current[276]), .y0(y0_current[276]));
  individual_277 dut_277(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[277]), .y2(y2_current[277]), .y1(y1_current[277]), .y0(y0_current[277]));
  individual_278 dut_278(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[278]), .y2(y2_current[278]), .y1(y1_current[278]), .y0(y0_current[278]));
  individual_279 dut_279(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[279]), .y2(y2_current[279]), .y1(y1_current[279]), .y0(y0_current[279]));
  individual_280 dut_280(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[280]), .y2(y2_current[280]), .y1(y1_current[280]), .y0(y0_current[280]));
  individual_281 dut_281(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[281]), .y2(y2_current[281]), .y1(y1_current[281]), .y0(y0_current[281]));
  individual_282 dut_282(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[282]), .y2(y2_current[282]), .y1(y1_current[282]), .y0(y0_current[282]));
  individual_283 dut_283(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[283]), .y2(y2_current[283]), .y1(y1_current[283]), .y0(y0_current[283]));
  individual_284 dut_284(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[284]), .y2(y2_current[284]), .y1(y1_current[284]), .y0(y0_current[284]));
  individual_285 dut_285(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[285]), .y2(y2_current[285]), .y1(y1_current[285]), .y0(y0_current[285]));
  individual_286 dut_286(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[286]), .y2(y2_current[286]), .y1(y1_current[286]), .y0(y0_current[286]));
  individual_287 dut_287(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[287]), .y2(y2_current[287]), .y1(y1_current[287]), .y0(y0_current[287]));
  individual_288 dut_288(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[288]), .y2(y2_current[288]), .y1(y1_current[288]), .y0(y0_current[288]));
  individual_289 dut_289(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[289]), .y2(y2_current[289]), .y1(y1_current[289]), .y0(y0_current[289]));
  individual_290 dut_290(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[290]), .y2(y2_current[290]), .y1(y1_current[290]), .y0(y0_current[290]));
  individual_291 dut_291(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[291]), .y2(y2_current[291]), .y1(y1_current[291]), .y0(y0_current[291]));
  individual_292 dut_292(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[292]), .y2(y2_current[292]), .y1(y1_current[292]), .y0(y0_current[292]));
  individual_293 dut_293(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[293]), .y2(y2_current[293]), .y1(y1_current[293]), .y0(y0_current[293]));
  individual_294 dut_294(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[294]), .y2(y2_current[294]), .y1(y1_current[294]), .y0(y0_current[294]));
  individual_295 dut_295(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[295]), .y2(y2_current[295]), .y1(y1_current[295]), .y0(y0_current[295]));
  individual_296 dut_296(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[296]), .y2(y2_current[296]), .y1(y1_current[296]), .y0(y0_current[296]));
  individual_297 dut_297(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[297]), .y2(y2_current[297]), .y1(y1_current[297]), .y0(y0_current[297]));
  individual_298 dut_298(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[298]), .y2(y2_current[298]), .y1(y1_current[298]), .y0(y0_current[298]));
  individual_299 dut_299(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[299]), .y2(y2_current[299]), .y1(y1_current[299]), .y0(y0_current[299]));
  individual_300 dut_300(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[300]), .y2(y2_current[300]), .y1(y1_current[300]), .y0(y0_current[300]));
  individual_301 dut_301(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[301]), .y2(y2_current[301]), .y1(y1_current[301]), .y0(y0_current[301]));
  individual_302 dut_302(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[302]), .y2(y2_current[302]), .y1(y1_current[302]), .y0(y0_current[302]));
  individual_303 dut_303(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[303]), .y2(y2_current[303]), .y1(y1_current[303]), .y0(y0_current[303]));
  individual_304 dut_304(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[304]), .y2(y2_current[304]), .y1(y1_current[304]), .y0(y0_current[304]));
  individual_305 dut_305(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[305]), .y2(y2_current[305]), .y1(y1_current[305]), .y0(y0_current[305]));
  individual_306 dut_306(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[306]), .y2(y2_current[306]), .y1(y1_current[306]), .y0(y0_current[306]));
  individual_307 dut_307(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[307]), .y2(y2_current[307]), .y1(y1_current[307]), .y0(y0_current[307]));
  individual_308 dut_308(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[308]), .y2(y2_current[308]), .y1(y1_current[308]), .y0(y0_current[308]));
  individual_309 dut_309(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[309]), .y2(y2_current[309]), .y1(y1_current[309]), .y0(y0_current[309]));
  individual_310 dut_310(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[310]), .y2(y2_current[310]), .y1(y1_current[310]), .y0(y0_current[310]));
  individual_311 dut_311(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[311]), .y2(y2_current[311]), .y1(y1_current[311]), .y0(y0_current[311]));
  individual_312 dut_312(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[312]), .y2(y2_current[312]), .y1(y1_current[312]), .y0(y0_current[312]));
  individual_313 dut_313(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[313]), .y2(y2_current[313]), .y1(y1_current[313]), .y0(y0_current[313]));
  individual_314 dut_314(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[314]), .y2(y2_current[314]), .y1(y1_current[314]), .y0(y0_current[314]));
  individual_315 dut_315(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[315]), .y2(y2_current[315]), .y1(y1_current[315]), .y0(y0_current[315]));
  individual_316 dut_316(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[316]), .y2(y2_current[316]), .y1(y1_current[316]), .y0(y0_current[316]));
  individual_317 dut_317(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[317]), .y2(y2_current[317]), .y1(y1_current[317]), .y0(y0_current[317]));
  individual_318 dut_318(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[318]), .y2(y2_current[318]), .y1(y1_current[318]), .y0(y0_current[318]));
  individual_319 dut_319(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[319]), .y2(y2_current[319]), .y1(y1_current[319]), .y0(y0_current[319]));
  individual_320 dut_320(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[320]), .y2(y2_current[320]), .y1(y1_current[320]), .y0(y0_current[320]));
  individual_321 dut_321(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[321]), .y2(y2_current[321]), .y1(y1_current[321]), .y0(y0_current[321]));
  individual_322 dut_322(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[322]), .y2(y2_current[322]), .y1(y1_current[322]), .y0(y0_current[322]));
  individual_323 dut_323(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[323]), .y2(y2_current[323]), .y1(y1_current[323]), .y0(y0_current[323]));
  individual_324 dut_324(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[324]), .y2(y2_current[324]), .y1(y1_current[324]), .y0(y0_current[324]));
  individual_325 dut_325(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[325]), .y2(y2_current[325]), .y1(y1_current[325]), .y0(y0_current[325]));
  individual_326 dut_326(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[326]), .y2(y2_current[326]), .y1(y1_current[326]), .y0(y0_current[326]));
  individual_327 dut_327(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[327]), .y2(y2_current[327]), .y1(y1_current[327]), .y0(y0_current[327]));
  individual_328 dut_328(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[328]), .y2(y2_current[328]), .y1(y1_current[328]), .y0(y0_current[328]));
  individual_329 dut_329(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[329]), .y2(y2_current[329]), .y1(y1_current[329]), .y0(y0_current[329]));
  individual_330 dut_330(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[330]), .y2(y2_current[330]), .y1(y1_current[330]), .y0(y0_current[330]));
  individual_331 dut_331(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[331]), .y2(y2_current[331]), .y1(y1_current[331]), .y0(y0_current[331]));
  individual_332 dut_332(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[332]), .y2(y2_current[332]), .y1(y1_current[332]), .y0(y0_current[332]));
  individual_333 dut_333(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[333]), .y2(y2_current[333]), .y1(y1_current[333]), .y0(y0_current[333]));
  individual_334 dut_334(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[334]), .y2(y2_current[334]), .y1(y1_current[334]), .y0(y0_current[334]));
  individual_335 dut_335(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[335]), .y2(y2_current[335]), .y1(y1_current[335]), .y0(y0_current[335]));
  individual_336 dut_336(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[336]), .y2(y2_current[336]), .y1(y1_current[336]), .y0(y0_current[336]));
  individual_337 dut_337(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[337]), .y2(y2_current[337]), .y1(y1_current[337]), .y0(y0_current[337]));
  individual_338 dut_338(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[338]), .y2(y2_current[338]), .y1(y1_current[338]), .y0(y0_current[338]));
  individual_339 dut_339(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[339]), .y2(y2_current[339]), .y1(y1_current[339]), .y0(y0_current[339]));
  individual_340 dut_340(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[340]), .y2(y2_current[340]), .y1(y1_current[340]), .y0(y0_current[340]));
  individual_341 dut_341(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[341]), .y2(y2_current[341]), .y1(y1_current[341]), .y0(y0_current[341]));
  individual_342 dut_342(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[342]), .y2(y2_current[342]), .y1(y1_current[342]), .y0(y0_current[342]));
  individual_343 dut_343(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[343]), .y2(y2_current[343]), .y1(y1_current[343]), .y0(y0_current[343]));
  individual_344 dut_344(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[344]), .y2(y2_current[344]), .y1(y1_current[344]), .y0(y0_current[344]));
  individual_345 dut_345(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[345]), .y2(y2_current[345]), .y1(y1_current[345]), .y0(y0_current[345]));
  individual_346 dut_346(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[346]), .y2(y2_current[346]), .y1(y1_current[346]), .y0(y0_current[346]));
  individual_347 dut_347(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[347]), .y2(y2_current[347]), .y1(y1_current[347]), .y0(y0_current[347]));
  individual_348 dut_348(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[348]), .y2(y2_current[348]), .y1(y1_current[348]), .y0(y0_current[348]));
  individual_349 dut_349(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[349]), .y2(y2_current[349]), .y1(y1_current[349]), .y0(y0_current[349]));
  individual_350 dut_350(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[350]), .y2(y2_current[350]), .y1(y1_current[350]), .y0(y0_current[350]));
  individual_351 dut_351(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[351]), .y2(y2_current[351]), .y1(y1_current[351]), .y0(y0_current[351]));
  individual_352 dut_352(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[352]), .y2(y2_current[352]), .y1(y1_current[352]), .y0(y0_current[352]));
  individual_353 dut_353(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[353]), .y2(y2_current[353]), .y1(y1_current[353]), .y0(y0_current[353]));
  individual_354 dut_354(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[354]), .y2(y2_current[354]), .y1(y1_current[354]), .y0(y0_current[354]));
  individual_355 dut_355(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[355]), .y2(y2_current[355]), .y1(y1_current[355]), .y0(y0_current[355]));
  individual_356 dut_356(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[356]), .y2(y2_current[356]), .y1(y1_current[356]), .y0(y0_current[356]));
  individual_357 dut_357(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[357]), .y2(y2_current[357]), .y1(y1_current[357]), .y0(y0_current[357]));
  individual_358 dut_358(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[358]), .y2(y2_current[358]), .y1(y1_current[358]), .y0(y0_current[358]));
  individual_359 dut_359(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[359]), .y2(y2_current[359]), .y1(y1_current[359]), .y0(y0_current[359]));
  individual_360 dut_360(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[360]), .y2(y2_current[360]), .y1(y1_current[360]), .y0(y0_current[360]));
  individual_361 dut_361(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[361]), .y2(y2_current[361]), .y1(y1_current[361]), .y0(y0_current[361]));
  individual_362 dut_362(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[362]), .y2(y2_current[362]), .y1(y1_current[362]), .y0(y0_current[362]));
  individual_363 dut_363(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[363]), .y2(y2_current[363]), .y1(y1_current[363]), .y0(y0_current[363]));
  individual_364 dut_364(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[364]), .y2(y2_current[364]), .y1(y1_current[364]), .y0(y0_current[364]));
  individual_365 dut_365(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[365]), .y2(y2_current[365]), .y1(y1_current[365]), .y0(y0_current[365]));
  individual_366 dut_366(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[366]), .y2(y2_current[366]), .y1(y1_current[366]), .y0(y0_current[366]));
  individual_367 dut_367(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[367]), .y2(y2_current[367]), .y1(y1_current[367]), .y0(y0_current[367]));
  individual_368 dut_368(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[368]), .y2(y2_current[368]), .y1(y1_current[368]), .y0(y0_current[368]));
  individual_369 dut_369(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[369]), .y2(y2_current[369]), .y1(y1_current[369]), .y0(y0_current[369]));
  individual_370 dut_370(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[370]), .y2(y2_current[370]), .y1(y1_current[370]), .y0(y0_current[370]));
  individual_371 dut_371(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[371]), .y2(y2_current[371]), .y1(y1_current[371]), .y0(y0_current[371]));
  individual_372 dut_372(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[372]), .y2(y2_current[372]), .y1(y1_current[372]), .y0(y0_current[372]));
  individual_373 dut_373(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[373]), .y2(y2_current[373]), .y1(y1_current[373]), .y0(y0_current[373]));
  individual_374 dut_374(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[374]), .y2(y2_current[374]), .y1(y1_current[374]), .y0(y0_current[374]));
  individual_375 dut_375(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[375]), .y2(y2_current[375]), .y1(y1_current[375]), .y0(y0_current[375]));
  individual_376 dut_376(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[376]), .y2(y2_current[376]), .y1(y1_current[376]), .y0(y0_current[376]));
  individual_377 dut_377(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[377]), .y2(y2_current[377]), .y1(y1_current[377]), .y0(y0_current[377]));
  individual_378 dut_378(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[378]), .y2(y2_current[378]), .y1(y1_current[378]), .y0(y0_current[378]));
  individual_379 dut_379(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[379]), .y2(y2_current[379]), .y1(y1_current[379]), .y0(y0_current[379]));
  individual_380 dut_380(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[380]), .y2(y2_current[380]), .y1(y1_current[380]), .y0(y0_current[380]));
  individual_381 dut_381(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[381]), .y2(y2_current[381]), .y1(y1_current[381]), .y0(y0_current[381]));
  individual_382 dut_382(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[382]), .y2(y2_current[382]), .y1(y1_current[382]), .y0(y0_current[382]));
  individual_383 dut_383(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[383]), .y2(y2_current[383]), .y1(y1_current[383]), .y0(y0_current[383]));
  individual_384 dut_384(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[384]), .y2(y2_current[384]), .y1(y1_current[384]), .y0(y0_current[384]));
  individual_385 dut_385(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[385]), .y2(y2_current[385]), .y1(y1_current[385]), .y0(y0_current[385]));
  individual_386 dut_386(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[386]), .y2(y2_current[386]), .y1(y1_current[386]), .y0(y0_current[386]));
  individual_387 dut_387(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[387]), .y2(y2_current[387]), .y1(y1_current[387]), .y0(y0_current[387]));
  individual_388 dut_388(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[388]), .y2(y2_current[388]), .y1(y1_current[388]), .y0(y0_current[388]));
  individual_389 dut_389(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[389]), .y2(y2_current[389]), .y1(y1_current[389]), .y0(y0_current[389]));
  individual_390 dut_390(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[390]), .y2(y2_current[390]), .y1(y1_current[390]), .y0(y0_current[390]));
  individual_391 dut_391(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[391]), .y2(y2_current[391]), .y1(y1_current[391]), .y0(y0_current[391]));
  individual_392 dut_392(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[392]), .y2(y2_current[392]), .y1(y1_current[392]), .y0(y0_current[392]));
  individual_393 dut_393(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[393]), .y2(y2_current[393]), .y1(y1_current[393]), .y0(y0_current[393]));
  individual_394 dut_394(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[394]), .y2(y2_current[394]), .y1(y1_current[394]), .y0(y0_current[394]));
  individual_395 dut_395(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[395]), .y2(y2_current[395]), .y1(y1_current[395]), .y0(y0_current[395]));
  individual_396 dut_396(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[396]), .y2(y2_current[396]), .y1(y1_current[396]), .y0(y0_current[396]));
  individual_397 dut_397(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[397]), .y2(y2_current[397]), .y1(y1_current[397]), .y0(y0_current[397]));
  individual_398 dut_398(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[398]), .y2(y2_current[398]), .y1(y1_current[398]), .y0(y0_current[398]));
  individual_399 dut_399(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[399]), .y2(y2_current[399]), .y1(y1_current[399]), .y0(y0_current[399]));
  individual_400 dut_400(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[400]), .y2(y2_current[400]), .y1(y1_current[400]), .y0(y0_current[400]));
  individual_401 dut_401(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[401]), .y2(y2_current[401]), .y1(y1_current[401]), .y0(y0_current[401]));
  individual_402 dut_402(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[402]), .y2(y2_current[402]), .y1(y1_current[402]), .y0(y0_current[402]));
  individual_403 dut_403(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[403]), .y2(y2_current[403]), .y1(y1_current[403]), .y0(y0_current[403]));
  individual_404 dut_404(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[404]), .y2(y2_current[404]), .y1(y1_current[404]), .y0(y0_current[404]));
  individual_405 dut_405(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[405]), .y2(y2_current[405]), .y1(y1_current[405]), .y0(y0_current[405]));
  individual_406 dut_406(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[406]), .y2(y2_current[406]), .y1(y1_current[406]), .y0(y0_current[406]));
  individual_407 dut_407(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[407]), .y2(y2_current[407]), .y1(y1_current[407]), .y0(y0_current[407]));
  individual_408 dut_408(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[408]), .y2(y2_current[408]), .y1(y1_current[408]), .y0(y0_current[408]));
  individual_409 dut_409(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[409]), .y2(y2_current[409]), .y1(y1_current[409]), .y0(y0_current[409]));
  individual_410 dut_410(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[410]), .y2(y2_current[410]), .y1(y1_current[410]), .y0(y0_current[410]));
  individual_411 dut_411(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[411]), .y2(y2_current[411]), .y1(y1_current[411]), .y0(y0_current[411]));
  individual_412 dut_412(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[412]), .y2(y2_current[412]), .y1(y1_current[412]), .y0(y0_current[412]));
  individual_413 dut_413(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[413]), .y2(y2_current[413]), .y1(y1_current[413]), .y0(y0_current[413]));
  individual_414 dut_414(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[414]), .y2(y2_current[414]), .y1(y1_current[414]), .y0(y0_current[414]));
  individual_415 dut_415(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[415]), .y2(y2_current[415]), .y1(y1_current[415]), .y0(y0_current[415]));
  individual_416 dut_416(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[416]), .y2(y2_current[416]), .y1(y1_current[416]), .y0(y0_current[416]));
  individual_417 dut_417(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[417]), .y2(y2_current[417]), .y1(y1_current[417]), .y0(y0_current[417]));
  individual_418 dut_418(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[418]), .y2(y2_current[418]), .y1(y1_current[418]), .y0(y0_current[418]));
  individual_419 dut_419(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[419]), .y2(y2_current[419]), .y1(y1_current[419]), .y0(y0_current[419]));
  individual_420 dut_420(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[420]), .y2(y2_current[420]), .y1(y1_current[420]), .y0(y0_current[420]));
  individual_421 dut_421(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[421]), .y2(y2_current[421]), .y1(y1_current[421]), .y0(y0_current[421]));
  individual_422 dut_422(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[422]), .y2(y2_current[422]), .y1(y1_current[422]), .y0(y0_current[422]));
  individual_423 dut_423(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[423]), .y2(y2_current[423]), .y1(y1_current[423]), .y0(y0_current[423]));
  individual_424 dut_424(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[424]), .y2(y2_current[424]), .y1(y1_current[424]), .y0(y0_current[424]));
  individual_425 dut_425(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[425]), .y2(y2_current[425]), .y1(y1_current[425]), .y0(y0_current[425]));
  individual_426 dut_426(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[426]), .y2(y2_current[426]), .y1(y1_current[426]), .y0(y0_current[426]));
  individual_427 dut_427(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[427]), .y2(y2_current[427]), .y1(y1_current[427]), .y0(y0_current[427]));
  individual_428 dut_428(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[428]), .y2(y2_current[428]), .y1(y1_current[428]), .y0(y0_current[428]));
  individual_429 dut_429(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[429]), .y2(y2_current[429]), .y1(y1_current[429]), .y0(y0_current[429]));
  individual_430 dut_430(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[430]), .y2(y2_current[430]), .y1(y1_current[430]), .y0(y0_current[430]));
  individual_431 dut_431(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[431]), .y2(y2_current[431]), .y1(y1_current[431]), .y0(y0_current[431]));
  individual_432 dut_432(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[432]), .y2(y2_current[432]), .y1(y1_current[432]), .y0(y0_current[432]));
  individual_433 dut_433(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[433]), .y2(y2_current[433]), .y1(y1_current[433]), .y0(y0_current[433]));
  individual_434 dut_434(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[434]), .y2(y2_current[434]), .y1(y1_current[434]), .y0(y0_current[434]));
  individual_435 dut_435(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[435]), .y2(y2_current[435]), .y1(y1_current[435]), .y0(y0_current[435]));
  individual_436 dut_436(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[436]), .y2(y2_current[436]), .y1(y1_current[436]), .y0(y0_current[436]));
  individual_437 dut_437(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[437]), .y2(y2_current[437]), .y1(y1_current[437]), .y0(y0_current[437]));
  individual_438 dut_438(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[438]), .y2(y2_current[438]), .y1(y1_current[438]), .y0(y0_current[438]));
  individual_439 dut_439(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[439]), .y2(y2_current[439]), .y1(y1_current[439]), .y0(y0_current[439]));
  individual_440 dut_440(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[440]), .y2(y2_current[440]), .y1(y1_current[440]), .y0(y0_current[440]));
  individual_441 dut_441(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[441]), .y2(y2_current[441]), .y1(y1_current[441]), .y0(y0_current[441]));
  individual_442 dut_442(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[442]), .y2(y2_current[442]), .y1(y1_current[442]), .y0(y0_current[442]));
  individual_443 dut_443(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[443]), .y2(y2_current[443]), .y1(y1_current[443]), .y0(y0_current[443]));
  individual_444 dut_444(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[444]), .y2(y2_current[444]), .y1(y1_current[444]), .y0(y0_current[444]));
  individual_445 dut_445(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[445]), .y2(y2_current[445]), .y1(y1_current[445]), .y0(y0_current[445]));
  individual_446 dut_446(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[446]), .y2(y2_current[446]), .y1(y1_current[446]), .y0(y0_current[446]));
  individual_447 dut_447(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[447]), .y2(y2_current[447]), .y1(y1_current[447]), .y0(y0_current[447]));
  individual_448 dut_448(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[448]), .y2(y2_current[448]), .y1(y1_current[448]), .y0(y0_current[448]));
  individual_449 dut_449(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[449]), .y2(y2_current[449]), .y1(y1_current[449]), .y0(y0_current[449]));
  individual_450 dut_450(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[450]), .y2(y2_current[450]), .y1(y1_current[450]), .y0(y0_current[450]));
  individual_451 dut_451(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[451]), .y2(y2_current[451]), .y1(y1_current[451]), .y0(y0_current[451]));
  individual_452 dut_452(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[452]), .y2(y2_current[452]), .y1(y1_current[452]), .y0(y0_current[452]));
  individual_453 dut_453(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[453]), .y2(y2_current[453]), .y1(y1_current[453]), .y0(y0_current[453]));
  individual_454 dut_454(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[454]), .y2(y2_current[454]), .y1(y1_current[454]), .y0(y0_current[454]));
  individual_455 dut_455(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[455]), .y2(y2_current[455]), .y1(y1_current[455]), .y0(y0_current[455]));
  individual_456 dut_456(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[456]), .y2(y2_current[456]), .y1(y1_current[456]), .y0(y0_current[456]));
  individual_457 dut_457(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[457]), .y2(y2_current[457]), .y1(y1_current[457]), .y0(y0_current[457]));
  individual_458 dut_458(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[458]), .y2(y2_current[458]), .y1(y1_current[458]), .y0(y0_current[458]));
  individual_459 dut_459(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[459]), .y2(y2_current[459]), .y1(y1_current[459]), .y0(y0_current[459]));
  individual_460 dut_460(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[460]), .y2(y2_current[460]), .y1(y1_current[460]), .y0(y0_current[460]));
  individual_461 dut_461(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[461]), .y2(y2_current[461]), .y1(y1_current[461]), .y0(y0_current[461]));
  individual_462 dut_462(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[462]), .y2(y2_current[462]), .y1(y1_current[462]), .y0(y0_current[462]));
  individual_463 dut_463(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[463]), .y2(y2_current[463]), .y1(y1_current[463]), .y0(y0_current[463]));
  individual_464 dut_464(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[464]), .y2(y2_current[464]), .y1(y1_current[464]), .y0(y0_current[464]));
  individual_465 dut_465(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[465]), .y2(y2_current[465]), .y1(y1_current[465]), .y0(y0_current[465]));
  individual_466 dut_466(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[466]), .y2(y2_current[466]), .y1(y1_current[466]), .y0(y0_current[466]));
  individual_467 dut_467(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[467]), .y2(y2_current[467]), .y1(y1_current[467]), .y0(y0_current[467]));
  individual_468 dut_468(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[468]), .y2(y2_current[468]), .y1(y1_current[468]), .y0(y0_current[468]));
  individual_469 dut_469(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[469]), .y2(y2_current[469]), .y1(y1_current[469]), .y0(y0_current[469]));
  individual_470 dut_470(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[470]), .y2(y2_current[470]), .y1(y1_current[470]), .y0(y0_current[470]));
  individual_471 dut_471(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[471]), .y2(y2_current[471]), .y1(y1_current[471]), .y0(y0_current[471]));
  individual_472 dut_472(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[472]), .y2(y2_current[472]), .y1(y1_current[472]), .y0(y0_current[472]));
  individual_473 dut_473(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[473]), .y2(y2_current[473]), .y1(y1_current[473]), .y0(y0_current[473]));
  individual_474 dut_474(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[474]), .y2(y2_current[474]), .y1(y1_current[474]), .y0(y0_current[474]));
  individual_475 dut_475(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[475]), .y2(y2_current[475]), .y1(y1_current[475]), .y0(y0_current[475]));
  individual_476 dut_476(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[476]), .y2(y2_current[476]), .y1(y1_current[476]), .y0(y0_current[476]));
  individual_477 dut_477(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[477]), .y2(y2_current[477]), .y1(y1_current[477]), .y0(y0_current[477]));
  individual_478 dut_478(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[478]), .y2(y2_current[478]), .y1(y1_current[478]), .y0(y0_current[478]));
  individual_479 dut_479(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[479]), .y2(y2_current[479]), .y1(y1_current[479]), .y0(y0_current[479]));
  individual_480 dut_480(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[480]), .y2(y2_current[480]), .y1(y1_current[480]), .y0(y0_current[480]));
  individual_481 dut_481(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[481]), .y2(y2_current[481]), .y1(y1_current[481]), .y0(y0_current[481]));
  individual_482 dut_482(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[482]), .y2(y2_current[482]), .y1(y1_current[482]), .y0(y0_current[482]));
  individual_483 dut_483(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[483]), .y2(y2_current[483]), .y1(y1_current[483]), .y0(y0_current[483]));
  individual_484 dut_484(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[484]), .y2(y2_current[484]), .y1(y1_current[484]), .y0(y0_current[484]));
  individual_485 dut_485(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[485]), .y2(y2_current[485]), .y1(y1_current[485]), .y0(y0_current[485]));
  individual_486 dut_486(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[486]), .y2(y2_current[486]), .y1(y1_current[486]), .y0(y0_current[486]));
  individual_487 dut_487(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[487]), .y2(y2_current[487]), .y1(y1_current[487]), .y0(y0_current[487]));
  individual_488 dut_488(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[488]), .y2(y2_current[488]), .y1(y1_current[488]), .y0(y0_current[488]));
  individual_489 dut_489(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[489]), .y2(y2_current[489]), .y1(y1_current[489]), .y0(y0_current[489]));
  individual_490 dut_490(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[490]), .y2(y2_current[490]), .y1(y1_current[490]), .y0(y0_current[490]));
  individual_491 dut_491(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[491]), .y2(y2_current[491]), .y1(y1_current[491]), .y0(y0_current[491]));
  individual_492 dut_492(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[492]), .y2(y2_current[492]), .y1(y1_current[492]), .y0(y0_current[492]));
  individual_493 dut_493(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[493]), .y2(y2_current[493]), .y1(y1_current[493]), .y0(y0_current[493]));
  individual_494 dut_494(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[494]), .y2(y2_current[494]), .y1(y1_current[494]), .y0(y0_current[494]));
  individual_495 dut_495(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[495]), .y2(y2_current[495]), .y1(y1_current[495]), .y0(y0_current[495]));
  individual_496 dut_496(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[496]), .y2(y2_current[496]), .y1(y1_current[496]), .y0(y0_current[496]));
  individual_497 dut_497(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[497]), .y2(y2_current[497]), .y1(y1_current[497]), .y0(y0_current[497]));
  individual_498 dut_498(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[498]), .y2(y2_current[498]), .y1(y1_current[498]), .y0(y0_current[498]));
  individual_499 dut_499(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[499]), .y2(y2_current[499]), .y1(y1_current[499]), .y0(y0_current[499]));
  individual_500 dut_500(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[500]), .y2(y2_current[500]), .y1(y1_current[500]), .y0(y0_current[500]));
  individual_501 dut_501(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[501]), .y2(y2_current[501]), .y1(y1_current[501]), .y0(y0_current[501]));
  individual_502 dut_502(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[502]), .y2(y2_current[502]), .y1(y1_current[502]), .y0(y0_current[502]));
  individual_503 dut_503(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[503]), .y2(y2_current[503]), .y1(y1_current[503]), .y0(y0_current[503]));
  individual_504 dut_504(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[504]), .y2(y2_current[504]), .y1(y1_current[504]), .y0(y0_current[504]));
  individual_505 dut_505(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[505]), .y2(y2_current[505]), .y1(y1_current[505]), .y0(y0_current[505]));
  individual_506 dut_506(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[506]), .y2(y2_current[506]), .y1(y1_current[506]), .y0(y0_current[506]));
  individual_507 dut_507(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[507]), .y2(y2_current[507]), .y1(y1_current[507]), .y0(y0_current[507]));
  individual_508 dut_508(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[508]), .y2(y2_current[508]), .y1(y1_current[508]), .y0(y0_current[508]));
  individual_509 dut_509(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[509]), .y2(y2_current[509]), .y1(y1_current[509]), .y0(y0_current[509]));
  individual_510 dut_510(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[510]), .y2(y2_current[510]), .y1(y1_current[510]), .y0(y0_current[510]));
  individual_511 dut_511(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[511]), .y2(y2_current[511]), .y1(y1_current[511]), .y0(y0_current[511]));
  individual_512 dut_512(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[512]), .y2(y2_current[512]), .y1(y1_current[512]), .y0(y0_current[512]));
  individual_513 dut_513(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[513]), .y2(y2_current[513]), .y1(y1_current[513]), .y0(y0_current[513]));
  individual_514 dut_514(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[514]), .y2(y2_current[514]), .y1(y1_current[514]), .y0(y0_current[514]));
  individual_515 dut_515(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[515]), .y2(y2_current[515]), .y1(y1_current[515]), .y0(y0_current[515]));
  individual_516 dut_516(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[516]), .y2(y2_current[516]), .y1(y1_current[516]), .y0(y0_current[516]));
  individual_517 dut_517(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[517]), .y2(y2_current[517]), .y1(y1_current[517]), .y0(y0_current[517]));
  individual_518 dut_518(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[518]), .y2(y2_current[518]), .y1(y1_current[518]), .y0(y0_current[518]));
  individual_519 dut_519(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[519]), .y2(y2_current[519]), .y1(y1_current[519]), .y0(y0_current[519]));
  individual_520 dut_520(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[520]), .y2(y2_current[520]), .y1(y1_current[520]), .y0(y0_current[520]));
  individual_521 dut_521(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[521]), .y2(y2_current[521]), .y1(y1_current[521]), .y0(y0_current[521]));
  individual_522 dut_522(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[522]), .y2(y2_current[522]), .y1(y1_current[522]), .y0(y0_current[522]));
  individual_523 dut_523(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[523]), .y2(y2_current[523]), .y1(y1_current[523]), .y0(y0_current[523]));
  individual_524 dut_524(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[524]), .y2(y2_current[524]), .y1(y1_current[524]), .y0(y0_current[524]));
  individual_525 dut_525(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[525]), .y2(y2_current[525]), .y1(y1_current[525]), .y0(y0_current[525]));
  individual_526 dut_526(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[526]), .y2(y2_current[526]), .y1(y1_current[526]), .y0(y0_current[526]));
  individual_527 dut_527(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[527]), .y2(y2_current[527]), .y1(y1_current[527]), .y0(y0_current[527]));
  individual_528 dut_528(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[528]), .y2(y2_current[528]), .y1(y1_current[528]), .y0(y0_current[528]));
  individual_529 dut_529(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[529]), .y2(y2_current[529]), .y1(y1_current[529]), .y0(y0_current[529]));
  individual_530 dut_530(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[530]), .y2(y2_current[530]), .y1(y1_current[530]), .y0(y0_current[530]));
  individual_531 dut_531(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[531]), .y2(y2_current[531]), .y1(y1_current[531]), .y0(y0_current[531]));
  individual_532 dut_532(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[532]), .y2(y2_current[532]), .y1(y1_current[532]), .y0(y0_current[532]));
  individual_533 dut_533(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[533]), .y2(y2_current[533]), .y1(y1_current[533]), .y0(y0_current[533]));
  individual_534 dut_534(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[534]), .y2(y2_current[534]), .y1(y1_current[534]), .y0(y0_current[534]));
  individual_535 dut_535(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[535]), .y2(y2_current[535]), .y1(y1_current[535]), .y0(y0_current[535]));
  individual_536 dut_536(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[536]), .y2(y2_current[536]), .y1(y1_current[536]), .y0(y0_current[536]));
  individual_537 dut_537(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[537]), .y2(y2_current[537]), .y1(y1_current[537]), .y0(y0_current[537]));
  individual_538 dut_538(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[538]), .y2(y2_current[538]), .y1(y1_current[538]), .y0(y0_current[538]));
  individual_539 dut_539(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[539]), .y2(y2_current[539]), .y1(y1_current[539]), .y0(y0_current[539]));
  individual_540 dut_540(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[540]), .y2(y2_current[540]), .y1(y1_current[540]), .y0(y0_current[540]));
  individual_541 dut_541(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[541]), .y2(y2_current[541]), .y1(y1_current[541]), .y0(y0_current[541]));
  individual_542 dut_542(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[542]), .y2(y2_current[542]), .y1(y1_current[542]), .y0(y0_current[542]));
  individual_543 dut_543(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[543]), .y2(y2_current[543]), .y1(y1_current[543]), .y0(y0_current[543]));
  individual_544 dut_544(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[544]), .y2(y2_current[544]), .y1(y1_current[544]), .y0(y0_current[544]));
  individual_545 dut_545(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[545]), .y2(y2_current[545]), .y1(y1_current[545]), .y0(y0_current[545]));
  individual_546 dut_546(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[546]), .y2(y2_current[546]), .y1(y1_current[546]), .y0(y0_current[546]));
  individual_547 dut_547(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[547]), .y2(y2_current[547]), .y1(y1_current[547]), .y0(y0_current[547]));
  individual_548 dut_548(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[548]), .y2(y2_current[548]), .y1(y1_current[548]), .y0(y0_current[548]));
  individual_549 dut_549(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[549]), .y2(y2_current[549]), .y1(y1_current[549]), .y0(y0_current[549]));
  individual_550 dut_550(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[550]), .y2(y2_current[550]), .y1(y1_current[550]), .y0(y0_current[550]));
  individual_551 dut_551(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[551]), .y2(y2_current[551]), .y1(y1_current[551]), .y0(y0_current[551]));
  individual_552 dut_552(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[552]), .y2(y2_current[552]), .y1(y1_current[552]), .y0(y0_current[552]));
  individual_553 dut_553(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[553]), .y2(y2_current[553]), .y1(y1_current[553]), .y0(y0_current[553]));
  individual_554 dut_554(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[554]), .y2(y2_current[554]), .y1(y1_current[554]), .y0(y0_current[554]));
  individual_555 dut_555(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[555]), .y2(y2_current[555]), .y1(y1_current[555]), .y0(y0_current[555]));
  individual_556 dut_556(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[556]), .y2(y2_current[556]), .y1(y1_current[556]), .y0(y0_current[556]));
  individual_557 dut_557(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[557]), .y2(y2_current[557]), .y1(y1_current[557]), .y0(y0_current[557]));
  individual_558 dut_558(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[558]), .y2(y2_current[558]), .y1(y1_current[558]), .y0(y0_current[558]));
  individual_559 dut_559(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[559]), .y2(y2_current[559]), .y1(y1_current[559]), .y0(y0_current[559]));
  individual_560 dut_560(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[560]), .y2(y2_current[560]), .y1(y1_current[560]), .y0(y0_current[560]));
  individual_561 dut_561(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[561]), .y2(y2_current[561]), .y1(y1_current[561]), .y0(y0_current[561]));
  individual_562 dut_562(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[562]), .y2(y2_current[562]), .y1(y1_current[562]), .y0(y0_current[562]));
  individual_563 dut_563(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[563]), .y2(y2_current[563]), .y1(y1_current[563]), .y0(y0_current[563]));
  individual_564 dut_564(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[564]), .y2(y2_current[564]), .y1(y1_current[564]), .y0(y0_current[564]));
  individual_565 dut_565(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[565]), .y2(y2_current[565]), .y1(y1_current[565]), .y0(y0_current[565]));
  individual_566 dut_566(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[566]), .y2(y2_current[566]), .y1(y1_current[566]), .y0(y0_current[566]));
  individual_567 dut_567(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[567]), .y2(y2_current[567]), .y1(y1_current[567]), .y0(y0_current[567]));
  individual_568 dut_568(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[568]), .y2(y2_current[568]), .y1(y1_current[568]), .y0(y0_current[568]));
  individual_569 dut_569(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[569]), .y2(y2_current[569]), .y1(y1_current[569]), .y0(y0_current[569]));
  individual_570 dut_570(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[570]), .y2(y2_current[570]), .y1(y1_current[570]), .y0(y0_current[570]));
  individual_571 dut_571(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[571]), .y2(y2_current[571]), .y1(y1_current[571]), .y0(y0_current[571]));
  individual_572 dut_572(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[572]), .y2(y2_current[572]), .y1(y1_current[572]), .y0(y0_current[572]));
  individual_573 dut_573(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[573]), .y2(y2_current[573]), .y1(y1_current[573]), .y0(y0_current[573]));
  individual_574 dut_574(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[574]), .y2(y2_current[574]), .y1(y1_current[574]), .y0(y0_current[574]));
  individual_575 dut_575(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[575]), .y2(y2_current[575]), .y1(y1_current[575]), .y0(y0_current[575]));
  individual_576 dut_576(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[576]), .y2(y2_current[576]), .y1(y1_current[576]), .y0(y0_current[576]));
  individual_577 dut_577(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[577]), .y2(y2_current[577]), .y1(y1_current[577]), .y0(y0_current[577]));
  individual_578 dut_578(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[578]), .y2(y2_current[578]), .y1(y1_current[578]), .y0(y0_current[578]));
  individual_579 dut_579(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[579]), .y2(y2_current[579]), .y1(y1_current[579]), .y0(y0_current[579]));
  individual_580 dut_580(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[580]), .y2(y2_current[580]), .y1(y1_current[580]), .y0(y0_current[580]));
  individual_581 dut_581(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[581]), .y2(y2_current[581]), .y1(y1_current[581]), .y0(y0_current[581]));
  individual_582 dut_582(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[582]), .y2(y2_current[582]), .y1(y1_current[582]), .y0(y0_current[582]));
  individual_583 dut_583(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[583]), .y2(y2_current[583]), .y1(y1_current[583]), .y0(y0_current[583]));
  individual_584 dut_584(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[584]), .y2(y2_current[584]), .y1(y1_current[584]), .y0(y0_current[584]));
  individual_585 dut_585(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[585]), .y2(y2_current[585]), .y1(y1_current[585]), .y0(y0_current[585]));
  individual_586 dut_586(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[586]), .y2(y2_current[586]), .y1(y1_current[586]), .y0(y0_current[586]));
  individual_587 dut_587(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[587]), .y2(y2_current[587]), .y1(y1_current[587]), .y0(y0_current[587]));
  individual_588 dut_588(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[588]), .y2(y2_current[588]), .y1(y1_current[588]), .y0(y0_current[588]));
  individual_589 dut_589(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[589]), .y2(y2_current[589]), .y1(y1_current[589]), .y0(y0_current[589]));
  individual_590 dut_590(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[590]), .y2(y2_current[590]), .y1(y1_current[590]), .y0(y0_current[590]));
  individual_591 dut_591(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[591]), .y2(y2_current[591]), .y1(y1_current[591]), .y0(y0_current[591]));
  individual_592 dut_592(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[592]), .y2(y2_current[592]), .y1(y1_current[592]), .y0(y0_current[592]));
  individual_593 dut_593(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[593]), .y2(y2_current[593]), .y1(y1_current[593]), .y0(y0_current[593]));
  individual_594 dut_594(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[594]), .y2(y2_current[594]), .y1(y1_current[594]), .y0(y0_current[594]));
  individual_595 dut_595(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[595]), .y2(y2_current[595]), .y1(y1_current[595]), .y0(y0_current[595]));
  individual_596 dut_596(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[596]), .y2(y2_current[596]), .y1(y1_current[596]), .y0(y0_current[596]));
  individual_597 dut_597(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[597]), .y2(y2_current[597]), .y1(y1_current[597]), .y0(y0_current[597]));
  individual_598 dut_598(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[598]), .y2(y2_current[598]), .y1(y1_current[598]), .y0(y0_current[598]));
  individual_599 dut_599(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[599]), .y2(y2_current[599]), .y1(y1_current[599]), .y0(y0_current[599]));
  individual_600 dut_600(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[600]), .y2(y2_current[600]), .y1(y1_current[600]), .y0(y0_current[600]));
  individual_601 dut_601(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[601]), .y2(y2_current[601]), .y1(y1_current[601]), .y0(y0_current[601]));
  individual_602 dut_602(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[602]), .y2(y2_current[602]), .y1(y1_current[602]), .y0(y0_current[602]));
  individual_603 dut_603(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[603]), .y2(y2_current[603]), .y1(y1_current[603]), .y0(y0_current[603]));
  individual_604 dut_604(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[604]), .y2(y2_current[604]), .y1(y1_current[604]), .y0(y0_current[604]));
  individual_605 dut_605(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[605]), .y2(y2_current[605]), .y1(y1_current[605]), .y0(y0_current[605]));
  individual_606 dut_606(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[606]), .y2(y2_current[606]), .y1(y1_current[606]), .y0(y0_current[606]));
  individual_607 dut_607(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[607]), .y2(y2_current[607]), .y1(y1_current[607]), .y0(y0_current[607]));
  individual_608 dut_608(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[608]), .y2(y2_current[608]), .y1(y1_current[608]), .y0(y0_current[608]));
  individual_609 dut_609(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[609]), .y2(y2_current[609]), .y1(y1_current[609]), .y0(y0_current[609]));
  individual_610 dut_610(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[610]), .y2(y2_current[610]), .y1(y1_current[610]), .y0(y0_current[610]));
  individual_611 dut_611(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[611]), .y2(y2_current[611]), .y1(y1_current[611]), .y0(y0_current[611]));
  individual_612 dut_612(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[612]), .y2(y2_current[612]), .y1(y1_current[612]), .y0(y0_current[612]));
  individual_613 dut_613(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[613]), .y2(y2_current[613]), .y1(y1_current[613]), .y0(y0_current[613]));
  individual_614 dut_614(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[614]), .y2(y2_current[614]), .y1(y1_current[614]), .y0(y0_current[614]));
  individual_615 dut_615(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[615]), .y2(y2_current[615]), .y1(y1_current[615]), .y0(y0_current[615]));
  individual_616 dut_616(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[616]), .y2(y2_current[616]), .y1(y1_current[616]), .y0(y0_current[616]));
  individual_617 dut_617(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[617]), .y2(y2_current[617]), .y1(y1_current[617]), .y0(y0_current[617]));
  individual_618 dut_618(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[618]), .y2(y2_current[618]), .y1(y1_current[618]), .y0(y0_current[618]));
  individual_619 dut_619(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[619]), .y2(y2_current[619]), .y1(y1_current[619]), .y0(y0_current[619]));
  individual_620 dut_620(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[620]), .y2(y2_current[620]), .y1(y1_current[620]), .y0(y0_current[620]));
  individual_621 dut_621(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[621]), .y2(y2_current[621]), .y1(y1_current[621]), .y0(y0_current[621]));
  individual_622 dut_622(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[622]), .y2(y2_current[622]), .y1(y1_current[622]), .y0(y0_current[622]));
  individual_623 dut_623(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[623]), .y2(y2_current[623]), .y1(y1_current[623]), .y0(y0_current[623]));
  individual_624 dut_624(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[624]), .y2(y2_current[624]), .y1(y1_current[624]), .y0(y0_current[624]));
  individual_625 dut_625(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[625]), .y2(y2_current[625]), .y1(y1_current[625]), .y0(y0_current[625]));
  individual_626 dut_626(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[626]), .y2(y2_current[626]), .y1(y1_current[626]), .y0(y0_current[626]));
  individual_627 dut_627(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[627]), .y2(y2_current[627]), .y1(y1_current[627]), .y0(y0_current[627]));
  individual_628 dut_628(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[628]), .y2(y2_current[628]), .y1(y1_current[628]), .y0(y0_current[628]));
  individual_629 dut_629(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[629]), .y2(y2_current[629]), .y1(y1_current[629]), .y0(y0_current[629]));
  individual_630 dut_630(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[630]), .y2(y2_current[630]), .y1(y1_current[630]), .y0(y0_current[630]));
  individual_631 dut_631(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[631]), .y2(y2_current[631]), .y1(y1_current[631]), .y0(y0_current[631]));
  individual_632 dut_632(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[632]), .y2(y2_current[632]), .y1(y1_current[632]), .y0(y0_current[632]));
  individual_633 dut_633(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[633]), .y2(y2_current[633]), .y1(y1_current[633]), .y0(y0_current[633]));
  individual_634 dut_634(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[634]), .y2(y2_current[634]), .y1(y1_current[634]), .y0(y0_current[634]));
  individual_635 dut_635(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[635]), .y2(y2_current[635]), .y1(y1_current[635]), .y0(y0_current[635]));
  individual_636 dut_636(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[636]), .y2(y2_current[636]), .y1(y1_current[636]), .y0(y0_current[636]));
  individual_637 dut_637(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[637]), .y2(y2_current[637]), .y1(y1_current[637]), .y0(y0_current[637]));
  individual_638 dut_638(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[638]), .y2(y2_current[638]), .y1(y1_current[638]), .y0(y0_current[638]));
  individual_639 dut_639(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[639]), .y2(y2_current[639]), .y1(y1_current[639]), .y0(y0_current[639]));
  individual_640 dut_640(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[640]), .y2(y2_current[640]), .y1(y1_current[640]), .y0(y0_current[640]));
  individual_641 dut_641(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[641]), .y2(y2_current[641]), .y1(y1_current[641]), .y0(y0_current[641]));
  individual_642 dut_642(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[642]), .y2(y2_current[642]), .y1(y1_current[642]), .y0(y0_current[642]));
  individual_643 dut_643(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[643]), .y2(y2_current[643]), .y1(y1_current[643]), .y0(y0_current[643]));
  individual_644 dut_644(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[644]), .y2(y2_current[644]), .y1(y1_current[644]), .y0(y0_current[644]));
  individual_645 dut_645(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[645]), .y2(y2_current[645]), .y1(y1_current[645]), .y0(y0_current[645]));
  individual_646 dut_646(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[646]), .y2(y2_current[646]), .y1(y1_current[646]), .y0(y0_current[646]));
  individual_647 dut_647(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[647]), .y2(y2_current[647]), .y1(y1_current[647]), .y0(y0_current[647]));
  individual_648 dut_648(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[648]), .y2(y2_current[648]), .y1(y1_current[648]), .y0(y0_current[648]));
  individual_649 dut_649(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[649]), .y2(y2_current[649]), .y1(y1_current[649]), .y0(y0_current[649]));
  individual_650 dut_650(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[650]), .y2(y2_current[650]), .y1(y1_current[650]), .y0(y0_current[650]));
  individual_651 dut_651(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[651]), .y2(y2_current[651]), .y1(y1_current[651]), .y0(y0_current[651]));
  individual_652 dut_652(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[652]), .y2(y2_current[652]), .y1(y1_current[652]), .y0(y0_current[652]));
  individual_653 dut_653(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[653]), .y2(y2_current[653]), .y1(y1_current[653]), .y0(y0_current[653]));
  individual_654 dut_654(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[654]), .y2(y2_current[654]), .y1(y1_current[654]), .y0(y0_current[654]));
  individual_655 dut_655(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[655]), .y2(y2_current[655]), .y1(y1_current[655]), .y0(y0_current[655]));
  individual_656 dut_656(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[656]), .y2(y2_current[656]), .y1(y1_current[656]), .y0(y0_current[656]));
  individual_657 dut_657(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[657]), .y2(y2_current[657]), .y1(y1_current[657]), .y0(y0_current[657]));
  individual_658 dut_658(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[658]), .y2(y2_current[658]), .y1(y1_current[658]), .y0(y0_current[658]));
  individual_659 dut_659(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[659]), .y2(y2_current[659]), .y1(y1_current[659]), .y0(y0_current[659]));
  individual_660 dut_660(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[660]), .y2(y2_current[660]), .y1(y1_current[660]), .y0(y0_current[660]));
  individual_661 dut_661(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[661]), .y2(y2_current[661]), .y1(y1_current[661]), .y0(y0_current[661]));
  individual_662 dut_662(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[662]), .y2(y2_current[662]), .y1(y1_current[662]), .y0(y0_current[662]));
  individual_663 dut_663(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[663]), .y2(y2_current[663]), .y1(y1_current[663]), .y0(y0_current[663]));
  individual_664 dut_664(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[664]), .y2(y2_current[664]), .y1(y1_current[664]), .y0(y0_current[664]));
  individual_665 dut_665(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[665]), .y2(y2_current[665]), .y1(y1_current[665]), .y0(y0_current[665]));
  individual_666 dut_666(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[666]), .y2(y2_current[666]), .y1(y1_current[666]), .y0(y0_current[666]));
  individual_667 dut_667(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[667]), .y2(y2_current[667]), .y1(y1_current[667]), .y0(y0_current[667]));
  individual_668 dut_668(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[668]), .y2(y2_current[668]), .y1(y1_current[668]), .y0(y0_current[668]));
  individual_669 dut_669(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[669]), .y2(y2_current[669]), .y1(y1_current[669]), .y0(y0_current[669]));
  individual_670 dut_670(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[670]), .y2(y2_current[670]), .y1(y1_current[670]), .y0(y0_current[670]));
  individual_671 dut_671(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[671]), .y2(y2_current[671]), .y1(y1_current[671]), .y0(y0_current[671]));
  individual_672 dut_672(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[672]), .y2(y2_current[672]), .y1(y1_current[672]), .y0(y0_current[672]));
  individual_673 dut_673(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[673]), .y2(y2_current[673]), .y1(y1_current[673]), .y0(y0_current[673]));
  individual_674 dut_674(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[674]), .y2(y2_current[674]), .y1(y1_current[674]), .y0(y0_current[674]));
  individual_675 dut_675(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[675]), .y2(y2_current[675]), .y1(y1_current[675]), .y0(y0_current[675]));
  individual_676 dut_676(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[676]), .y2(y2_current[676]), .y1(y1_current[676]), .y0(y0_current[676]));
  individual_677 dut_677(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[677]), .y2(y2_current[677]), .y1(y1_current[677]), .y0(y0_current[677]));
  individual_678 dut_678(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[678]), .y2(y2_current[678]), .y1(y1_current[678]), .y0(y0_current[678]));
  individual_679 dut_679(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[679]), .y2(y2_current[679]), .y1(y1_current[679]), .y0(y0_current[679]));
  individual_680 dut_680(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[680]), .y2(y2_current[680]), .y1(y1_current[680]), .y0(y0_current[680]));
  individual_681 dut_681(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[681]), .y2(y2_current[681]), .y1(y1_current[681]), .y0(y0_current[681]));
  individual_682 dut_682(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[682]), .y2(y2_current[682]), .y1(y1_current[682]), .y0(y0_current[682]));
  individual_683 dut_683(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[683]), .y2(y2_current[683]), .y1(y1_current[683]), .y0(y0_current[683]));
  individual_684 dut_684(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[684]), .y2(y2_current[684]), .y1(y1_current[684]), .y0(y0_current[684]));
  individual_685 dut_685(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[685]), .y2(y2_current[685]), .y1(y1_current[685]), .y0(y0_current[685]));
  individual_686 dut_686(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[686]), .y2(y2_current[686]), .y1(y1_current[686]), .y0(y0_current[686]));
  individual_687 dut_687(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[687]), .y2(y2_current[687]), .y1(y1_current[687]), .y0(y0_current[687]));
  individual_688 dut_688(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[688]), .y2(y2_current[688]), .y1(y1_current[688]), .y0(y0_current[688]));
  individual_689 dut_689(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[689]), .y2(y2_current[689]), .y1(y1_current[689]), .y0(y0_current[689]));
  individual_690 dut_690(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[690]), .y2(y2_current[690]), .y1(y1_current[690]), .y0(y0_current[690]));
  individual_691 dut_691(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[691]), .y2(y2_current[691]), .y1(y1_current[691]), .y0(y0_current[691]));
  individual_692 dut_692(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[692]), .y2(y2_current[692]), .y1(y1_current[692]), .y0(y0_current[692]));
  individual_693 dut_693(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[693]), .y2(y2_current[693]), .y1(y1_current[693]), .y0(y0_current[693]));
  individual_694 dut_694(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[694]), .y2(y2_current[694]), .y1(y1_current[694]), .y0(y0_current[694]));
  individual_695 dut_695(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[695]), .y2(y2_current[695]), .y1(y1_current[695]), .y0(y0_current[695]));
  individual_696 dut_696(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[696]), .y2(y2_current[696]), .y1(y1_current[696]), .y0(y0_current[696]));
  individual_697 dut_697(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[697]), .y2(y2_current[697]), .y1(y1_current[697]), .y0(y0_current[697]));
  individual_698 dut_698(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[698]), .y2(y2_current[698]), .y1(y1_current[698]), .y0(y0_current[698]));
  individual_699 dut_699(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[699]), .y2(y2_current[699]), .y1(y1_current[699]), .y0(y0_current[699]));
  individual_700 dut_700(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[700]), .y2(y2_current[700]), .y1(y1_current[700]), .y0(y0_current[700]));
  individual_701 dut_701(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[701]), .y2(y2_current[701]), .y1(y1_current[701]), .y0(y0_current[701]));
  individual_702 dut_702(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[702]), .y2(y2_current[702]), .y1(y1_current[702]), .y0(y0_current[702]));
  individual_703 dut_703(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[703]), .y2(y2_current[703]), .y1(y1_current[703]), .y0(y0_current[703]));
  individual_704 dut_704(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[704]), .y2(y2_current[704]), .y1(y1_current[704]), .y0(y0_current[704]));
  individual_705 dut_705(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[705]), .y2(y2_current[705]), .y1(y1_current[705]), .y0(y0_current[705]));
  individual_706 dut_706(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[706]), .y2(y2_current[706]), .y1(y1_current[706]), .y0(y0_current[706]));
  individual_707 dut_707(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[707]), .y2(y2_current[707]), .y1(y1_current[707]), .y0(y0_current[707]));
  individual_708 dut_708(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[708]), .y2(y2_current[708]), .y1(y1_current[708]), .y0(y0_current[708]));
  individual_709 dut_709(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[709]), .y2(y2_current[709]), .y1(y1_current[709]), .y0(y0_current[709]));
  individual_710 dut_710(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[710]), .y2(y2_current[710]), .y1(y1_current[710]), .y0(y0_current[710]));
  individual_711 dut_711(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[711]), .y2(y2_current[711]), .y1(y1_current[711]), .y0(y0_current[711]));
  individual_712 dut_712(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[712]), .y2(y2_current[712]), .y1(y1_current[712]), .y0(y0_current[712]));
  individual_713 dut_713(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[713]), .y2(y2_current[713]), .y1(y1_current[713]), .y0(y0_current[713]));
  individual_714 dut_714(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[714]), .y2(y2_current[714]), .y1(y1_current[714]), .y0(y0_current[714]));
  individual_715 dut_715(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[715]), .y2(y2_current[715]), .y1(y1_current[715]), .y0(y0_current[715]));
  individual_716 dut_716(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[716]), .y2(y2_current[716]), .y1(y1_current[716]), .y0(y0_current[716]));
  individual_717 dut_717(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[717]), .y2(y2_current[717]), .y1(y1_current[717]), .y0(y0_current[717]));
  individual_718 dut_718(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[718]), .y2(y2_current[718]), .y1(y1_current[718]), .y0(y0_current[718]));
  individual_719 dut_719(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[719]), .y2(y2_current[719]), .y1(y1_current[719]), .y0(y0_current[719]));
  individual_720 dut_720(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[720]), .y2(y2_current[720]), .y1(y1_current[720]), .y0(y0_current[720]));
  individual_721 dut_721(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[721]), .y2(y2_current[721]), .y1(y1_current[721]), .y0(y0_current[721]));
  individual_722 dut_722(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[722]), .y2(y2_current[722]), .y1(y1_current[722]), .y0(y0_current[722]));
  individual_723 dut_723(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[723]), .y2(y2_current[723]), .y1(y1_current[723]), .y0(y0_current[723]));
  individual_724 dut_724(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[724]), .y2(y2_current[724]), .y1(y1_current[724]), .y0(y0_current[724]));
  individual_725 dut_725(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[725]), .y2(y2_current[725]), .y1(y1_current[725]), .y0(y0_current[725]));
  individual_726 dut_726(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[726]), .y2(y2_current[726]), .y1(y1_current[726]), .y0(y0_current[726]));
  individual_727 dut_727(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[727]), .y2(y2_current[727]), .y1(y1_current[727]), .y0(y0_current[727]));
  individual_728 dut_728(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[728]), .y2(y2_current[728]), .y1(y1_current[728]), .y0(y0_current[728]));
  individual_729 dut_729(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[729]), .y2(y2_current[729]), .y1(y1_current[729]), .y0(y0_current[729]));
  individual_730 dut_730(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[730]), .y2(y2_current[730]), .y1(y1_current[730]), .y0(y0_current[730]));
  individual_731 dut_731(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[731]), .y2(y2_current[731]), .y1(y1_current[731]), .y0(y0_current[731]));
  individual_732 dut_732(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[732]), .y2(y2_current[732]), .y1(y1_current[732]), .y0(y0_current[732]));
  individual_733 dut_733(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[733]), .y2(y2_current[733]), .y1(y1_current[733]), .y0(y0_current[733]));
  individual_734 dut_734(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[734]), .y2(y2_current[734]), .y1(y1_current[734]), .y0(y0_current[734]));
  individual_735 dut_735(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[735]), .y2(y2_current[735]), .y1(y1_current[735]), .y0(y0_current[735]));
  individual_736 dut_736(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[736]), .y2(y2_current[736]), .y1(y1_current[736]), .y0(y0_current[736]));
  individual_737 dut_737(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[737]), .y2(y2_current[737]), .y1(y1_current[737]), .y0(y0_current[737]));
  individual_738 dut_738(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[738]), .y2(y2_current[738]), .y1(y1_current[738]), .y0(y0_current[738]));
  individual_739 dut_739(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[739]), .y2(y2_current[739]), .y1(y1_current[739]), .y0(y0_current[739]));
  individual_740 dut_740(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[740]), .y2(y2_current[740]), .y1(y1_current[740]), .y0(y0_current[740]));
  individual_741 dut_741(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[741]), .y2(y2_current[741]), .y1(y1_current[741]), .y0(y0_current[741]));
  individual_742 dut_742(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[742]), .y2(y2_current[742]), .y1(y1_current[742]), .y0(y0_current[742]));
  individual_743 dut_743(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[743]), .y2(y2_current[743]), .y1(y1_current[743]), .y0(y0_current[743]));
  individual_744 dut_744(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[744]), .y2(y2_current[744]), .y1(y1_current[744]), .y0(y0_current[744]));
  individual_745 dut_745(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[745]), .y2(y2_current[745]), .y1(y1_current[745]), .y0(y0_current[745]));
  individual_746 dut_746(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[746]), .y2(y2_current[746]), .y1(y1_current[746]), .y0(y0_current[746]));
  individual_747 dut_747(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[747]), .y2(y2_current[747]), .y1(y1_current[747]), .y0(y0_current[747]));
  individual_748 dut_748(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[748]), .y2(y2_current[748]), .y1(y1_current[748]), .y0(y0_current[748]));
  individual_749 dut_749(.a1(a1), .a0(a0), .b1(b1), .b0(b0), .y3(y3_current[749]), .y2(y2_current[749]), .y1(y1_current[749]), .y0(y0_current[749]));

	// Create task to evaluate each testcase
	// Note that this evaluates the entire population for this testcase
	task testcase;
		input [15:0] a1_value;
input [15:0] a0_value;
input [15:0] b1_value;
input [15:0] b0_value;
input [15:0] y3_value;
input [15:0] y2_value;
input [15:0] y1_value;
input [15:0] y0_value;


		// Initialise inputs
		a1=a1_value;
		a0=a0_value;
		b1=b1_value;
		b0=b0_value;

		for(int i = 0; i < `POPULATION_SIZE; i++) begin
 // calculate hamming distance
 fitness[i]  = $countones(~(y3_current[i]  ^ y3_value)) + $countones(~(y2_current[i]  ^ y2_value)) + $countones(~(y1_current[i]  ^ y1_value)) + $countones(~(y0_current[i]  ^ y0_value));

		end
	endtask

	// We want to change our inputs on negedge so that we can run testcases at posedge
	always @(posedge clk) begin
		if (rst == 0) begin
			{a1, a0, b1, b0, y3_expected, y2_expected, y1_expected, y0_expected} = testvectors[vectornum];
			vectornum = vectornum + 1;
			testcase(a1, a0, b1, b0, y3_expected, y2_expected, y1_expected, y0_expected);
		end

	if (vectornum == `TEST_COUNT) begin
		// Print all fitness scores to the console
		for(int i = 0; i < `POPULATION_SIZE; i++) begin
			$display("%0d",fitness[i]);
		end

		$stop;

	end

end

  // We use a clock to load in our testvectors
  always begin
    #(`PERIOD/2) clk = ~clk;
  end

  // Run simulation
  initial begin
  
    // Set all scores to zero
    for(int i = 0; i < `POPULATION_SIZE; i++) begin
      fitness[i] = 0;
    end
       
    // Set the clock high so we get posedges at 10,20,30 etc.
    //clk = 1;
    clk = 1; rst = 1;
    #(`PERIOD) rst = 0;

    // DEBUGGING - Dump to vcd file
    //$dumpfile("testbench_values.vcd");
    //$dumpvars(0,fulladder_tb);

    // Read in test vectors
    $readmemb("template/test_vectors.tv", testvectors);
    // test vectors
    //$writememb("tmp/memory_b.txt",testvectors);
	
    
    // Wait clock cycles for test to complete
    #(`PERIOD*`TEST_COUNT);
    
    // Print all fitness scores to the console
    //for(int i = 0; i < `POPULATION_SIZE; i++) begin
      //$display("%0d",fitness[i]);
    //end

    $finish;
  end
 endmodule
