input logic clock
input logic reset
input logic i
output logic out
