
      endcase
    end
  end
endmodule
