input wire clk
input wire rst
input wire j
input wire k
output reg q
