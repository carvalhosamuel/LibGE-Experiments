module mux(output logic out, input logic a0, a1, a2, d0, d1, d2, d3, d4, d5, d6, d7);
  always@(*) begin
