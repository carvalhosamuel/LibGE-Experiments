input logic [15:0] a1
input logic [15:0] a0
input logic [15:0] b1
input logic [15:0] b0
output logic [15:0] y3
output logic [15:0] y2
output logic [15:0] y1
output logic [15:0] y0
