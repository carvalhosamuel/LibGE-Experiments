input wire clk
input wire rst
input wire sel
output reg [2:0] q
