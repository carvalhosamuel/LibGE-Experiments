      if(q_current[i] == q_value) begin
          fitness[i] = fitness[i] + 1;
      end
