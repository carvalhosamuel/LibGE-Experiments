input wire a
input wire b
input wire ci
output wire sum
output wire co
