module ssd(output logic[6:0] seg, input logic[3:0] bcd);
  always @(*) begin
