
  
endmodule
