  end
endmodule
